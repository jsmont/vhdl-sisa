library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity font_rom is
    generic (data_width  : natural := 8;
             addr_length : natural := 12);
    port (clk :in std_logic;
          address :in std_logic_vector(addr_length-1 downto 0);
          data_out:out std_logic_vector(data_width-1 downto 0));
end font_rom;

architecture synth of font_rom is

	constant mem_size : natural := 2**addr_length;
	type mem_type is array (mem_size-1 downto 0) of std_logic_vector (data_width-1 downto 0);

	constant mem : mem_type := (
-- 0x00 ''
0=> "01111110",      --   ****** 
1=> "11000011",      --  **    **
2=> "10011001",      --  *  **  *
3=> "10011001",      --  *  **  *
4=> "11110011",      --  ****  **
5=> "11100111",      --  ***  ***
6=> "11100111",      --  ***  ***
7=> "11111111",      --  ********
8=> "11100111",      --  ***  ***
9=> "11100111",      --  ***  ***
10=> "01111110",     --   ****** 
11=> "00000000",     --          
-- 0x01 ''         
12=> "00000000",     --          
13=> "00000000",     --          
14=> "00000000",     --          
15=> "01110110",     --   *** ** 
16=> "11011100",     --  ** ***  
17=> "00000000",     --          
18=> "01110110",     --   *** ** 
19=> "11011100",     --  ** ***  
20=> "00000000",     --          
21=> "00000000",     --          
22=> "00000000",     --          
23=> "00000000",     --          
-- 0x02 ''         
24=> "01101110",     --   ** *** 
25=> "11011000",     --  ** **   
26=> "11011000",     --  ** **   
27=> "11011000",     --  ** **   
28=> "11011000",     --  ** **   
29=> "11011110",     --  ** **** 
30=> "11011000",     --  ** **   
31=> "11011000",     --  ** **   
32=> "11011000",     --  ** **   
33=> "01101110",     --   ** *** 
34=> "00000000",     --          
35=> "00000000",     --          
-- 0x03 ''         
36=> "00000000",     --          
37=> "00000000",     --          
38=> "00000000",     --          
39=> "01101110",     --   ** *** 
40=> "11011011",     --  ** ** **
41=> "11011011",     --  ** ** **
42=> "11011111",     --  ** *****
43=> "11011000",     --  ** **   
44=> "11011011",     --  ** ** **
45=> "01101110",     --   ** *** 
46=> "00000000",     --          
47=> "00000000",     --          
-- 0x04 ''         
48=> "00000000",     --          
49=> "00000000",     --          
50=> "00010000",     --     *    
51=> "00111000",     --    ***   
52=> "01111100",     --   *****  
53=> "11111110",     --  ******* 
54=> "01111100",     --   *****  
55=> "00111000",     --    ***   
56=> "00010000",     --     *    
57=> "00000000",     --          
58=> "00000000",     --          
59=> "00000000",     --          
-- 0x05 ''         
60=> "10001000",     --  *   *   
61=> "10001000",     --  *   *   
62=> "11111000",     --  *****   
63=> "10001000",     --  *   *   
64=> "10001000",     --  *   *   
65=> "00000000",     --          
66=> "00111110",     --    ***** 
67=> "00001000",     --      *   
68=> "00001000",     --      *   
69=> "00001000",     --      *   
70=> "00001000",     --      *   
71=> "00000000",     --          
-- 0x06 ''         
72=> "11111000",     --  *****   
73=> "10000000",     --  *       
74=> "11100000",     --  ***     
75=> "10000000",     --  *       
76=> "10000000",     --  *       
77=> "00000000",     --          
78=> "00111110",     --    ***** 
79=> "00100000",     --    *     
80=> "00111000",     --    ***   
81=> "00100000",     --    *     
82=> "00100000",     --    *     
83=> "00000000",     --          
-- 0x07 ''         
84=> "01111000",     --   ****   
85=> "10000000",     --  *       
86=> "10000000",     --  *       
87=> "10000000",     --  *       
88=> "01111000",     --   ****   
89=> "00000000",     --          
90=> "00111100",     --    ****  
91=> "00100010",     --    *   * 
92=> "00111110",     --    ***** 
93=> "00100100",     --    *  *  
94=> "00100010",     --    *   * 
95=> "00000000",     --          
-- 0x08 ''         
96=> "10000000",     --  *       
97=> "10000000",     --  *       
98=> "10000000",     --  *       
99=> "10000000",     --  *       
100=> "11111000",    --  *****   
101=> "00000000",    --          
102=> "00111110",    --    ***** 
103=> "00100000",    --    *     
104=> "00111000",    --    ***   
105=> "00100000",    --    *     
106=> "00100000",    --    *     
107=> "00000000",    --          
-- 0x09 ''         
108=> "00100010",    --    *   * 
109=> "10001000",    --  *   *   
110=> "00100010",    --    *   * 
111=> "10001000",    --  *   *   
112=> "00100010",    --    *   * 
113=> "10001000",    --  *   *   
114=> "00100010",    --    *   * 
115=> "10001000",    --  *   *   
116=> "00100010",    --    *   * 
117=> "10001000",    --  *   *   
118=> "00100010",    --    *   * 
119=> "10001000",    --  *   *   
-- 0x0A ''         
120=> "01010101",    --   * * * *
121=> "10101010",    --  * * * * 
122=> "01010101",    --   * * * *
123=> "10101010",    --  * * * * 
124=> "01010101",    --   * * * *
125=> "10101010",    --  * * * * 
126=> "01010101",    --   * * * *
127=> "10101010",    --  * * * * 
128=> "01010101",    --   * * * *
129=> "10101010",    --  * * * * 
130=> "01010101",    --   * * * *
131=> "10101010",    --  * * * * 
-- 0x0B ''         
132=> "11101110",    --  *** *** 
133=> "10111011",    --  * *** **
134=> "11101110",    --  *** *** 
135=> "10111011",    --  * *** **
136=> "11101110",    --  *** *** 
137=> "10111011",    --  * *** **
138=> "11101110",    --  *** *** 
139=> "10111011",    --  * *** **
140=> "11101110",    --  *** *** 
141=> "10111011",    --  * *** **
142=> "11101110",    --  *** *** 
143=> "10111011",    --  * *** **
-- 0x0C ''         
144=> "11111111",    --  ********
145=> "11111111",    --  ********
146=> "11111111",    --  ********
147=> "11111111",    --  ********
148=> "11111111",    --  ********
149=> "11111111",    --  ********
150=> "11111111",    --  ********
151=> "11111111",    --  ********
152=> "11111111",    --  ********
153=> "11111111",    --  ********
154=> "11111111",    --  ********
155=> "11111111",    --  ********
-- 0x0D ''         
156=> "00000000",    --          
157=> "00000000",    --          
158=> "00000000",    --          
159=> "00000000",    --          
160=> "00000000",    --          
161=> "00000000",    --          
162=> "11111111",    --  ********
163=> "11111111",    --  ********
164=> "11111111",    --  ********
165=> "11111111",    --  ********
166=> "11111111",    --  ********
167=> "11111111",    --  ********
-- 0x0E ''         
168=> "11111111",    --  ********
169=> "11111111",    --  ********
170=> "11111111",    --  ********
171=> "11111111",    --  ********
172=> "11111111",    --  ********
173=> "11111111",    --  ********
174=> "00000000",    --          
175=> "00000000",    --          
176=> "00000000",    --          
177=> "00000000",    --          
178=> "00000000",    --          
179=> "00000000",    --          
-- 0x0F ''         
180=> "11110000",    --  ****    
181=> "11110000",    --  ****    
182=> "11110000",    --  ****    
183=> "11110000",    --  ****    
184=> "11110000",    --  ****    
185=> "11110000",    --  ****    
186=> "11110000",    --  ****    
187=> "11110000",    --  ****    
188=> "11110000",    --  ****    
189=> "11110000",    --  ****    
190=> "11110000",    --  ****    
191=> "11110000",    --  ****    
-- 0x10 ''         
192=> "00001111",    --      ****
193=> "00001111",    --      ****
194=> "00001111",    --      ****
195=> "00001111",    --      ****
196=> "00001111",    --      ****
197=> "00001111",    --      ****
198=> "00001111",    --      ****
199=> "00001111",    --      ****
200=> "00001111",    --      ****
201=> "00001111",    --      ****
202=> "00001111",    --      ****
203=> "00001111",    --      ****
-- 0x11 ''         
204=> "10001000",    --  *   *   
205=> "11001000",    --  **  *   
206=> "10101000",    --  * * *   
207=> "10011000",    --  *  **   
208=> "10001000",    --  *   *   
209=> "00000000",    --          
210=> "00100000",    --    *     
211=> "00100000",    --    *     
212=> "00100000",    --    *     
213=> "00100000",    --    *     
214=> "00111110",    --    ***** 
215=> "00000000",    --          
-- 0x12 ''         
216=> "10001000",    --  *   *   
217=> "10001000",    --  *   *   
218=> "01010000",    --   * *    
219=> "01010000",    --   * *    
220=> "00100000",    --    *     
221=> "00000000",    --          
222=> "00111110",    --    ***** 
223=> "00001000",    --      *   
224=> "00001000",    --      *   
225=> "00001000",    --      *   
226=> "00001000",    --      *   
227=> "00000000",    --          
-- 0x13 ''         
228=> "00000000",    --          
229=> "00000000",    --          
230=> "00000110",    --       ** 
231=> "00001100",    --      **  
232=> "00011000",    --     **   
233=> "00110000",    --    **    
234=> "01111110",    --   ****** 
235=> "00000000",    --          
236=> "01111110",    --   ****** 
237=> "00000000",    --          
238=> "00000000",    --          
239=> "00000000",    --          
-- 0x14 ''         
240=> "00000000",    --          
241=> "00000000",    --          
242=> "01100000",    --   **     
243=> "00110000",    --    **    
244=> "00011000",    --     **   
245=> "00001100",    --      **  
246=> "01111110",    --   ****** 
247=> "00000000",    --          
248=> "01111110",    --   ****** 
249=> "00000000",    --          
250=> "00000000",    --          
251=> "00000000",    --          
-- 0x15 ''         
252=> "00000000",    --          
253=> "00000000",    --          
254=> "00000110",    --       ** 
255=> "00001100",    --      **  
256=> "11111110",    --  ******* 
257=> "00111000",    --    ***   
258=> "11111110",    --  ******* 
259=> "01100000",    --   **     
260=> "11000000",    --  **      
261=> "00000000",    --          
262=> "00000000",    --          
263=> "00000000",    --          
-- 0x16 ''         
264=> "00000000",    --          
265=> "00000010",    --        * 
266=> "00001110",    --      *** 
267=> "00111110",    --    ***** 
268=> "01111110",    --   ****** 
269=> "11111110",    --  ******* 
270=> "01111110",    --   ****** 
271=> "00111110",    --    ***** 
272=> "00001110",    --      *** 
273=> "00000010",    --        * 
274=> "00000000",    --          
275=> "00000000",    --          
-- 0x17 ''         
276=> "00000000",    --          
277=> "10000000",    --  *       
278=> "11100000",    --  ***     
279=> "11110000",    --  ****    
280=> "11111100",    --  ******  
281=> "11111110",    --  ******* 
282=> "11111100",    --  ******  
283=> "11110000",    --  ****    
284=> "11100000",    --  ***     
285=> "10000000",    --  *       
286=> "00000000",    --          
287=> "00000000",    --          
-- 0x18 ''         
288=> "00000000",    --          
289=> "00011000",    --     **   
290=> "00111100",    --    ****  
291=> "01111110",    --   ****** 
292=> "00011000",    --     **   
293=> "00011000",    --     **   
294=> "00011000",    --     **   
295=> "00011000",    --     **   
296=> "00011000",    --     **   
297=> "00011000",    --     **   
298=> "00000000",    --          
299=> "00000000",    --          
-- 0x19 ''         
300=> "00000000",    --          
301=> "00011000",    --     **   
302=> "00011000",    --     **   
303=> "00011000",    --     **   
304=> "00011000",    --     **   
305=> "00011000",    --     **   
306=> "00011000",    --     **   
307=> "01111110",    --   ****** 
308=> "00111100",    --    ****  
309=> "00011000",    --     **   
310=> "00000000",    --          
311=> "00000000",    --          
-- 0x1A ''         
312=> "00000000",    --          
313=> "00000000",    --          
314=> "00000000",    --          
315=> "00011000",    --     **   
316=> "00001100",    --      **  
317=> "11111110",    --  ******* 
318=> "00001100",    --      **  
319=> "00011000",    --     **   
320=> "00000000",    --          
321=> "00000000",    --          
322=> "00000000",    --          
323=> "00000000",    --          
-- 0x1B ''         
324=> "00000000",    --          
325=> "00000000",    --          
326=> "00000000",    --          
327=> "00110000",    --    **    
328=> "01100000",    --   **     
329=> "11111110",    --  ******* 
330=> "01100000",    --   **     
331=> "00110000",    --    **    
332=> "00000000",    --          
333=> "00000000",    --          
334=> "00000000",    --          
335=> "00000000",    --          
-- 0x1C ''         
336=> "00000000",    --          
337=> "00011000",    --     **   
338=> "00111100",    --    ****  
339=> "01111110",    --   ****** 
340=> "00011000",    --     **   
341=> "00011000",    --     **   
342=> "00011000",    --     **   
343=> "01111110",    --   ****** 
344=> "00111100",    --    ****  
345=> "00011000",    --     **   
346=> "00000000",    --          
347=> "00000000",    --          
-- 0x1D ''         
348=> "00000000",    --          
349=> "00000000",    --          
350=> "00000000",    --          
351=> "00101000",    --    * *   
352=> "01101100",    --   ** **  
353=> "11111110",    --  ******* 
354=> "01101100",    --   ** **  
355=> "00101000",    --    * *   
356=> "00000000",    --          
357=> "00000000",    --          
358=> "00000000",    --          
359=> "00000000",    --          
-- 0x1E ''         
360=> "00000000",    --          
361=> "00000110",    --       ** 
362=> "00000110",    --       ** 
363=> "00110110",    --    ** ** 
364=> "01100110",    --   **  ** 
365=> "11111110",    --  ******* 
366=> "01100000",    --   **     
367=> "00110000",    --    **    
368=> "00000000",    --          
369=> "00000000",    --          
370=> "00000000",    --          
371=> "00000000",    --          
-- 0x1F ''         
372=> "00000000",    --          
373=> "00000000",    --          
374=> "00000000",    --          
375=> "11000000",    --  **      
376=> "01111100",    --   *****  
377=> "01101110",    --   ** *** 
378=> "01101100",    --   ** **  
379=> "01101100",    --   ** **  
380=> "01101100",    --   ** **  
381=> "00000000",    --          
382=> "00000000",    --          
383=> "00000000",    --          
-- 0x20 ' '        
384=> "00000000",    --          
385=> "00000000",    --          
386=> "00000000",    --          
387=> "00000000",    --          
388=> "00000000",    --          
389=> "00000000",    --          
390=> "00000000",    --          
391=> "00000000",    --          
392=> "00000000",    --          
393=> "00000000",    --          
394=> "00000000",    --          
395=> "00000000",    --          
-- 0x21 '!'        
396=> "00000000",    --          
397=> "00011000",    --     **   
398=> "00111100",    --    ****  
399=> "00111100",    --    ****  
400=> "00111100",    --    ****  
401=> "00011000",    --     **   
402=> "00011000",    --     **   
403=> "00000000",    --          
404=> "00011000",    --     **   
405=> "00011000",    --     **   
406=> "00000000",    --          
407=> "00000000",    --          
-- 0x22 '"'        
408=> "00000000",    --          
409=> "00110110",    --    ** ** 
410=> "00110110",    --    ** ** 
411=> "00010100",    --     * *  
412=> "00000000",    --          
413=> "00000000",    --          
414=> "00000000",    --          
415=> "00000000",    --          
416=> "00000000",    --          
417=> "00000000",    --          
418=> "00000000",    --          
419=> "00000000",    --          
-- 0x23 '#'        
420=> "00000000",    --          
421=> "00000000",    --          
422=> "00000000",    --          
423=> "01101100",    --   ** **  
424=> "11111110",    --  ******* 
425=> "01101100",    --   ** **  
426=> "01101100",    --   ** **  
427=> "01101100",    --   ** **  
428=> "11111110",    --  ******* 
429=> "01101100",    --   ** **  
430=> "00000000",    --          
431=> "00000000",    --          
-- 0x24 '$'        
432=> "00000000",    --          
433=> "00010000",    --     *    
434=> "01111100",    --   *****  
435=> "11010110",    --  ** * ** 
436=> "01110000",    --   ***    
437=> "00111000",    --    ***   
438=> "00011100",    --     ***  
439=> "11010110",    --  ** * ** 
440=> "01111100",    --   *****  
441=> "00010000",    --     *    
442=> "00000000",    --          
443=> "00000000",    --          
-- 0x25 '%'        
444=> "00000000",    --          
445=> "00000000",    --          
446=> "00000000",    --          
447=> "01100010",    --   **   * 
448=> "01100110",    --   **  ** 
449=> "00001100",    --      **  
450=> "00011000",    --     **   
451=> "00110000",    --    **    
452=> "01100110",    --   **  ** 
453=> "11000110",    --  **   ** 
454=> "00000000",    --          
455=> "00000000",    --          
-- 0x26 '&'        
456=> "00000000",    --          
457=> "00111000",    --    ***   
458=> "01101100",    --   ** **  
459=> "00111000",    --    ***   
460=> "00111000",    --    ***   
461=> "01110010",    --   ***  * 
462=> "11111110",    --  ******* 
463=> "11001100",    --  **  **  
464=> "11001100",    --  **  **  
465=> "01110110",    --   *** ** 
466=> "00000000",    --          
467=> "00000000",    --          
-- 0x27 "'"        
468=> "00011100",    --     ***  
469=> "00011100",    --     ***  
470=> "00001100",    --      **  
471=> "00011000",    --     **   
472=> "00000000",    --          
473=> "00000000",    --          
474=> "00000000",    --          
475=> "00000000",    --          
476=> "00000000",    --          
477=> "00000000",    --          
478=> "00000000",    --          
479=> "00000000",    --          
-- 0x28 '('        
480=> "00000000",    --          
481=> "00001100",    --      **  
482=> "00011000",    --     **   
483=> "00110000",    --    **    
484=> "00110000",    --    **    
485=> "00110000",    --    **    
486=> "00110000",    --    **    
487=> "00110000",    --    **    
488=> "00011000",    --     **   
489=> "00001100",    --      **  
490=> "00000000",    --          
491=> "00000000",    --          
-- 0x29 ')'        
492=> "00000000",    --          
493=> "00110000",    --    **    
494=> "00011000",    --     **   
495=> "00001100",    --      **  
496=> "00001100",    --      **  
497=> "00001100",    --      **  
498=> "00001100",    --      **  
499=> "00001100",    --      **  
500=> "00011000",    --     **   
501=> "00110000",    --    **    
502=> "00000000",    --          
503=> "00000000",    --          
-- 0x2A '*'        
504=> "00000000",    --          
505=> "00000000",    --          
506=> "00000000",    --          
507=> "01101100",    --   ** **  
508=> "00111000",    --    ***   
509=> "11111110",    --  ******* 
510=> "00111000",    --    ***   
511=> "01101100",    --   ** **  
512=> "00000000",    --          
513=> "00000000",    --          
514=> "00000000",    --          
515=> "00000000",    --          
-- 0x2B '+'        
516=> "00000000",    --          
517=> "00000000",    --          
518=> "00000000",    --          
519=> "00011000",    --     **   
520=> "00011000",    --     **   
521=> "01111110",    --   ****** 
522=> "00011000",    --     **   
523=> "00011000",    --     **   
524=> "00000000",    --          
525=> "00000000",    --          
526=> "00000000",    --          
527=> "00000000",    --          
-- 0x2C ','        
528=> "00000000",    --          
529=> "00000000",    --          
530=> "00000000",    --          
531=> "00000000",    --          
532=> "00000000",    --          
533=> "00000000",    --          
534=> "00000000",    --          
535=> "00001100",    --      **  
536=> "00001100",    --      **  
537=> "00001100",    --      **  
538=> "00011000",    --     **   
539=> "00000000",    --          
-- 0x2D '-'        
540=> "00000000",    --          
541=> "00000000",    --          
542=> "00000000",    --          
543=> "00000000",    --          
544=> "00000000",    --          
545=> "11111110",    --  ******* 
546=> "00000000",    --          
547=> "00000000",    --          
548=> "00000000",    --          
549=> "00000000",    --          
550=> "00000000",    --          
551=> "00000000",    --          
-- 0x2E '.'        
552=> "00000000",    --          
553=> "00000000",    --          
554=> "00000000",    --          
555=> "00000000",    --          
556=> "00000000",    --          
557=> "00000000",    --          
558=> "00000000",    --          
559=> "00000000",    --          
560=> "00011000",    --     **   
561=> "00011000",    --     **   
562=> "00000000",    --          
563=> "00000000",    --          
-- 0x2F '/'        
564=> "00000000",    --          
565=> "00000000",    --          
566=> "00000000",    --          
567=> "00000110",    --       ** 
568=> "00001100",    --      **  
569=> "00011000",    --     **   
570=> "00110000",    --    **    
571=> "01100000",    --   **     
572=> "11000000",    --  **      
573=> "00000000",    --          
574=> "00000000",    --          
575=> "00000000",    --          
-- 0x30 '0'        
576=> "00000000",    --          
577=> "01111100",    --   *****  
578=> "11000110",    --  **   ** 
579=> "11000110",    --  **   ** 
580=> "11000110",    --  **   ** 
581=> "11010110",    --  ** * ** 
582=> "11000110",    --  **   ** 
583=> "11000110",    --  **   ** 
584=> "11000110",    --  **   ** 
585=> "01111100",    --   *****  
586=> "00000000",    --          
587=> "00000000",    --          
-- 0x31 '1'        
588=> "00000000",    --          
589=> "00011000",    --     **   
590=> "01111000",    --   ****   
591=> "00011000",    --     **   
592=> "00011000",    --     **   
593=> "00011000",    --     **   
594=> "00011000",    --     **   
595=> "00011000",    --     **   
596=> "00011000",    --     **   
597=> "01111110",    --   ****** 
598=> "00000000",    --          
599=> "00000000",    --          
-- 0x32 '2'        
600=> "00000000",    --          
601=> "01111100",    --   *****  
602=> "11000110",    --  **   ** 
603=> "11000110",    --  **   ** 
604=> "00001100",    --      **  
605=> "00011000",    --     **   
606=> "00110000",    --    **    
607=> "01100000",    --   **     
608=> "11000110",    --  **   ** 
609=> "11111110",    --  ******* 
610=> "00000000",    --          
611=> "00000000",    --          
-- 0x33 '3'        
612=> "00000000",    --          
613=> "01111100",    --   *****  
614=> "11000110",    --  **   ** 
615=> "00000110",    --       ** 
616=> "00000110",    --       ** 
617=> "00111100",    --    ****  
618=> "00000110",    --       ** 
619=> "00000110",    --       ** 
620=> "11000110",    --  **   ** 
621=> "01111100",    --   *****  
622=> "00000000",    --          
623=> "00000000",    --          
-- 0x34 '4'        
624=> "00000000",    --          
625=> "00001100",    --      **  
626=> "00011100",    --     ***  
627=> "00111100",    --    ****  
628=> "01101100",    --   ** **  
629=> "11001100",    --  **  **  
630=> "11111110",    --  ******* 
631=> "00001100",    --      **  
632=> "00001100",    --      **  
633=> "00001100",    --      **  
634=> "00000000",    --          
635=> "00000000",    --          
-- 0x35 '5'        
636=> "00000000",    --          
637=> "11111110",    --  ******* 
638=> "11000000",    --  **      
639=> "11000000",    --  **      
640=> "11000000",    --  **      
641=> "11111100",    --  ******  
642=> "00000110",    --       ** 
643=> "00000110",    --       ** 
644=> "11000110",    --  **   ** 
645=> "01111100",    --   *****  
646=> "00000000",    --          
647=> "00000000",    --          
-- 0x36 '6'        
648=> "00000000",    --          
649=> "01111100",    --   *****  
650=> "11000110",    --  **   ** 
651=> "11000000",    --  **      
652=> "11000000",    --  **      
653=> "11111100",    --  ******  
654=> "11000110",    --  **   ** 
655=> "11000110",    --  **   ** 
656=> "11000110",    --  **   ** 
657=> "01111100",    --   *****  
658=> "00000000",    --          
659=> "00000000",    --          
-- 0x37 '7'        
660=> "00000000",    --          
661=> "11111110",    --  ******* 
662=> "11000110",    --  **   ** 
663=> "00001100",    --      **  
664=> "00011000",    --     **   
665=> "00110000",    --    **    
666=> "00110000",    --    **    
667=> "00110000",    --    **    
668=> "00110000",    --    **    
669=> "00110000",    --    **    
670=> "00000000",    --          
671=> "00000000",    --          
-- 0x38 '8'        
672=> "00000000",    --          
673=> "01111100",    --   *****  
674=> "11000110",    --  **   ** 
675=> "11000110",    --  **   ** 
676=> "11000110",    --  **   ** 
677=> "01111100",    --   *****  
678=> "11000110",    --  **   ** 
679=> "11000110",    --  **   ** 
680=> "11000110",    --  **   ** 
681=> "01111100",    --   *****  
682=> "00000000",    --          
683=> "00000000",    --          
-- 0x39 '9'        
684=> "00000000",    --          
685=> "01111100",    --   *****  
686=> "11000110",    --  **   ** 
687=> "11000110",    --  **   ** 
688=> "11000110",    --  **   ** 
689=> "01111110",    --   ****** 
690=> "00000110",    --       ** 
691=> "00000110",    --       ** 
692=> "11000110",    --  **   ** 
693=> "01111100",    --   *****  
694=> "00000000",    --          
695=> "00000000",    --          
-- 0x3A ':'        
696=> "00000000",    --          
697=> "00000000",    --          
698=> "00000000",    --          
699=> "00001100",    --      **  
700=> "00001100",    --      **  
701=> "00000000",    --          
702=> "00000000",    --          
703=> "00001100",    --      **  
704=> "00001100",    --      **  
705=> "00000000",    --          
706=> "00000000",    --          
707=> "00000000",    --          
-- 0x3B ';'        
708=> "00000000",    --          
709=> "00000000",    --          
710=> "00000000",    --          
711=> "00001100",    --      **  
712=> "00001100",    --      **  
713=> "00000000",    --          
714=> "00000000",    --          
715=> "00001100",    --      **  
716=> "00001100",    --      **  
717=> "00001100",    --      **  
718=> "00011000",    --     **   
719=> "00000000",    --          
-- 0x3C '<'        
720=> "00000000",    --          
721=> "00001100",    --      **  
722=> "00011000",    --     **   
723=> "00110000",    --    **    
724=> "01100000",    --   **     
725=> "11000000",    --  **      
726=> "01100000",    --   **     
727=> "00110000",    --    **    
728=> "00011000",    --     **   
729=> "00001100",    --      **  
730=> "00000000",    --          
731=> "00000000",    --          
-- 0x3D '='        
732=> "00000000",    --          
733=> "00000000",    --          
734=> "00000000",    --          
735=> "00000000",    --          
736=> "11111110",    --  ******* 
737=> "00000000",    --          
738=> "11111110",    --  ******* 
739=> "00000000",    --          
740=> "00000000",    --          
741=> "00000000",    --          
742=> "00000000",    --          
743=> "00000000",    --          
-- 0x3E '>'        
744=> "00000000",    --          
745=> "01100000",    --   **     
746=> "00110000",    --    **    
747=> "00011000",    --     **   
748=> "00001100",    --      **  
749=> "00000110",    --       ** 
750=> "00001100",    --      **  
751=> "00011000",    --     **   
752=> "00110000",    --    **    
753=> "01100000",    --   **     
754=> "00000000",    --          
755=> "00000000",    --          
-- 0x3F '?'        
756=> "00000000",    --          
757=> "01111100",    --   *****  
758=> "11000110",    --  **   ** 
759=> "11000110",    --  **   ** 
760=> "00001100",    --      **  
761=> "00011000",    --     **   
762=> "00011000",    --     **   
763=> "00000000",    --          
764=> "00011000",    --     **   
765=> "00011000",    --     **   
766=> "00000000",    --          
767=> "00000000",    --          
-- 0x40 '@'        
768=> "00000000",    --          
769=> "01111100",    --   *****  
770=> "11000110",    --  **   ** 
771=> "11000110",    --  **   ** 
772=> "11011110",    --  ** **** 
773=> "11011110",    --  ** **** 
774=> "11011110",    --  ** **** 
775=> "11011100",    --  ** ***  
776=> "11000000",    --  **      
777=> "01111110",    --   ****** 
778=> "00000000",    --          
779=> "00000000",    --          
-- 0x41 'A'        
780=> "00000000",    --          
781=> "00111000",    --    ***   
782=> "01101100",    --   ** **  
783=> "11000110",    --  **   ** 
784=> "11000110",    --  **   ** 
785=> "11000110",    --  **   ** 
786=> "11111110",    --  ******* 
787=> "11000110",    --  **   ** 
788=> "11000110",    --  **   ** 
789=> "11000110",    --  **   ** 
790=> "00000000",    --          
791=> "00000000",    --          
-- 0x42 'B'        
792=> "00000000",    --          
793=> "11111100",    --  ******  
794=> "01100110",    --   **  ** 
795=> "01100110",    --   **  ** 
796=> "01100110",    --   **  ** 
797=> "01111100",    --   *****  
798=> "01100110",    --   **  ** 
799=> "01100110",    --   **  ** 
800=> "01100110",    --   **  ** 
801=> "11111100",    --  ******  
802=> "00000000",    --          
803=> "00000000",    --          
-- 0x43 'C'        
804=> "00000000",    --          
805=> "00111100",    --    ****  
806=> "01100110",    --   **  ** 
807=> "11000000",    --  **      
808=> "11000000",    --  **      
809=> "11000000",    --  **      
810=> "11000000",    --  **      
811=> "11000000",    --  **      
812=> "01100110",    --   **  ** 
813=> "00111100",    --    ****  
814=> "00000000",    --          
815=> "00000000",    --          
-- 0x44 'D'        
816=> "00000000",    --          
817=> "11111000",    --  *****   
818=> "01101100",    --   ** **  
819=> "01100110",    --   **  ** 
820=> "01100110",    --   **  ** 
821=> "01100110",    --   **  ** 
822=> "01100110",    --   **  ** 
823=> "01100110",    --   **  ** 
824=> "01101100",    --   ** **  
825=> "11111000",    --  *****   
826=> "00000000",    --          
827=> "00000000",    --          
-- 0x45 'E'        
828=> "00000000",    --          
829=> "11111110",    --  ******* 
830=> "01100110",    --   **  ** 
831=> "01100000",    --   **     
832=> "01100000",    --   **     
833=> "01111100",    --   *****  
834=> "01100000",    --   **     
835=> "01100000",    --   **     
836=> "01100110",    --   **  ** 
837=> "11111110",    --  ******* 
838=> "00000000",    --          
839=> "00000000",    --          
-- 0x46 'F'        
840=> "00000000",    --          
841=> "11111110",    --  ******* 
842=> "01100110",    --   **  ** 
843=> "01100000",    --   **     
844=> "01100000",    --   **     
845=> "01111100",    --   *****  
846=> "01100000",    --   **     
847=> "01100000",    --   **     
848=> "01100000",    --   **     
849=> "11110000",    --  ****    
850=> "00000000",    --          
851=> "00000000",    --          
-- 0x47 'G'        
852=> "00000000",    --          
853=> "01111100",    --   *****  
854=> "11000110",    --  **   ** 
855=> "11000110",    --  **   ** 
856=> "11000000",    --  **      
857=> "11000000",    --  **      
858=> "11001110",    --  **  *** 
859=> "11000110",    --  **   ** 
860=> "11000110",    --  **   ** 
861=> "01111100",    --   *****  
862=> "00000000",    --          
863=> "00000000",    --          
-- 0x48 'H'        
864=> "00000000",    --          
865=> "11000110",    --  **   ** 
866=> "11000110",    --  **   ** 
867=> "11000110",    --  **   ** 
868=> "11000110",    --  **   ** 
869=> "11111110",    --  ******* 
870=> "11000110",    --  **   ** 
871=> "11000110",    --  **   ** 
872=> "11000110",    --  **   ** 
873=> "11000110",    --  **   ** 
874=> "00000000",    --          
875=> "00000000",    --          
-- 0x49 'I'        
876=> "00000000",    --          
877=> "00111100",    --    ****  
878=> "00011000",    --     **   
879=> "00011000",    --     **   
880=> "00011000",    --     **   
881=> "00011000",    --     **   
882=> "00011000",    --     **   
883=> "00011000",    --     **   
884=> "00011000",    --     **   
885=> "00111100",    --    ****  
886=> "00000000",    --          
887=> "00000000",    --          
-- 0x4A 'J'        
888=> "00000000",    --          
889=> "00111100",    --    ****  
890=> "00011000",    --     **   
891=> "00011000",    --     **   
892=> "00011000",    --     **   
893=> "00011000",    --     **   
894=> "00011000",    --     **   
895=> "11011000",    --  ** **   
896=> "11011000",    --  ** **   
897=> "01110000",    --   ***    
898=> "00000000",    --          
899=> "00000000",    --          
-- 0x4B 'K'        
900=> "00000000",    --          
901=> "11000110",    --  **   ** 
902=> "11001100",    --  **  **  
903=> "11011000",    --  ** **   
904=> "11110000",    --  ****    
905=> "11110000",    --  ****    
906=> "11011000",    --  ** **   
907=> "11001100",    --  **  **  
908=> "11000110",    --  **   ** 
909=> "11000110",    --  **   ** 
910=> "00000000",    --          
911=> "00000000",    --          
-- 0x4C 'L'        
912=> "00000000",    --          
913=> "11110000",    --  ****    
914=> "01100000",    --   **     
915=> "01100000",    --   **     
916=> "01100000",    --   **     
917=> "01100000",    --   **     
918=> "01100000",    --   **     
919=> "01100010",    --   **   * 
920=> "01100110",    --   **  ** 
921=> "11111110",    --  ******* 
922=> "00000000",    --          
923=> "00000000",    --          
-- 0x4D 'M'        
924=> "00000000",    --          
925=> "11000110",    --  **   ** 
926=> "11000110",    --  **   ** 
927=> "11101110",    --  *** *** 
928=> "11111110",    --  ******* 
929=> "11010110",    --  ** * ** 
930=> "11010110",    --  ** * ** 
931=> "11010110",    --  ** * ** 
932=> "11000110",    --  **   ** 
933=> "11000110",    --  **   ** 
934=> "00000000",    --          
935=> "00000000",    --          
-- 0x4E 'N'        
936=> "00000000",    --          
937=> "11000110",    --  **   ** 
938=> "11000110",    --  **   ** 
939=> "11100110",    --  ***  ** 
940=> "11100110",    --  ***  ** 
941=> "11110110",    --  **** ** 
942=> "11011110",    --  ** **** 
943=> "11001110",    --  **  *** 
944=> "11001110",    --  **  *** 
945=> "11000110",    --  **   ** 
946=> "00000000",    --          
947=> "00000000",    --          
-- 0x4F 'O'        
948=> "00000000",    --          
949=> "01111100",    --   *****  
950=> "11000110",    --  **   ** 
951=> "11000110",    --  **   ** 
952=> "11000110",    --  **   ** 
953=> "11000110",    --  **   ** 
954=> "11000110",    --  **   ** 
955=> "11000110",    --  **   ** 
956=> "11000110",    --  **   ** 
957=> "01111100",    --   *****  
958=> "00000000",    --          
959=> "00000000",    --          
-- 0x50 'P'        
960=> "00000000",    --          
961=> "11111100",    --  ******  
962=> "01100110",    --   **  ** 
963=> "01100110",    --   **  ** 
964=> "01100110",    --   **  ** 
965=> "01111100",    --   *****  
966=> "01100000",    --   **     
967=> "01100000",    --   **     
968=> "01100000",    --   **     
969=> "11110000",    --  ****    
970=> "00000000",    --          
971=> "00000000",    --          
-- 0x51 'Q'        
972=> "00000000",    --          
973=> "01111100",    --   *****  
974=> "11000110",    --  **   ** 
975=> "11000110",    --  **   ** 
976=> "11000110",    --  **   ** 
977=> "11000110",    --  **   ** 
978=> "11000110",    --  **   ** 
979=> "11000110",    --  **   ** 
980=> "11010110",    --  ** * ** 
981=> "01111100",    --   *****  
982=> "00000110",    --       ** 
983=> "00000000",    --          
-- 0x52 'R'        
984=> "00000000",    --          
985=> "11111100",    --  ******  
986=> "01100110",    --   **  ** 
987=> "01100110",    --   **  ** 
988=> "01100110",    --   **  ** 
989=> "01111100",    --   *****  
990=> "01111000",    --   ****   
991=> "01101100",    --   ** **  
992=> "01100110",    --   **  ** 
993=> "11100110",    --  ***  ** 
994=> "00000000",    --          
995=> "00000000",    --          
-- 0x53 'S'        
996=> "00000000",    --          
997=> "01111100",    --   *****  
998=> "11000110",    --  **   ** 
999=> "11000000",    --  **      
1000=> "01100000",   --   **     
1001=> "00111000",   --    ***   
1002=> "00001100",   --      **  
1003=> "00000110",   --       ** 
1004=> "11000110",   --  **   ** 
1005=> "01111100",   --   *****  
1006=> "00000000",   --          
1007=> "00000000",   --          
-- 0x54 'T'        
1008=> "00000000",   --          
1009=> "01111110",   --   ****** 
1010=> "01011010",   --   * ** * 
1011=> "00011000",   --     **   
1012=> "00011000",   --     **   
1013=> "00011000",   --     **   
1014=> "00011000",   --     **   
1015=> "00011000",   --     **   
1016=> "00011000",   --     **   
1017=> "00111100",   --    ****  
1018=> "00000000",   --          
1019=> "00000000",   --          
-- 0x55 'U'        
1020=> "00000000",   --          
1021=> "11000110",   --  **   ** 
1022=> "11000110",   --  **   ** 
1023=> "11000110",   --  **   ** 
1024=> "11000110",   --  **   ** 
1025=> "11000110",   --  **   ** 
1026=> "11000110",   --  **   ** 
1027=> "11000110",   --  **   ** 
1028=> "11000110",   --  **   ** 
1029=> "01111100",   --   *****  
1030=> "00000000",   --          
1031=> "00000000",   --          
-- 0x56 'V'        
1032=> "00000000",   --          
1033=> "11000110",   --  **   ** 
1034=> "11000110",   --  **   ** 
1035=> "11000110",   --  **   ** 
1036=> "11000110",   --  **   ** 
1037=> "11000110",   --  **   ** 
1038=> "11000110",   --  **   ** 
1039=> "01101100",   --   ** **  
1040=> "00111000",   --    ***   
1041=> "00010000",   --     *    
1042=> "00000000",   --          
1043=> "00000000",   --          
-- 0x57 'W'        
1044=> "00000000",   --          
1045=> "11000110",   --  **   ** 
1046=> "11000110",   --  **   ** 
1047=> "11010110",   --  ** * ** 
1048=> "11010110",   --  ** * ** 
1049=> "11010110",   --  ** * ** 
1050=> "11111110",   --  ******* 
1051=> "11101110",   --  *** *** 
1052=> "11000110",   --  **   ** 
1053=> "11000110",   --  **   ** 
1054=> "00000000",   --          
1055=> "00000000",   --          
-- 0x58 'X'        
1056=> "00000000",   --          
1057=> "11000110",   --  **   ** 
1058=> "11000110",   --  **   ** 
1059=> "01101100",   --   ** **  
1060=> "00111000",   --    ***   
1061=> "00111000",   --    ***   
1062=> "00111000",   --    ***   
1063=> "01101100",   --   ** **  
1064=> "11000110",   --  **   ** 
1065=> "11000110",   --  **   ** 
1066=> "00000000",   --          
1067=> "00000000",   --          
-- 0x59 'Y'        
1068=> "00000000",   --          
1069=> "01100110",   --   **  ** 
1070=> "01100110",   --   **  ** 
1071=> "01100110",   --   **  ** 
1072=> "01100110",   --   **  ** 
1073=> "00111100",   --    ****  
1074=> "00011000",   --     **   
1075=> "00011000",   --     **   
1076=> "00011000",   --     **   
1077=> "00111100",   --    ****  
1078=> "00000000",   --          
1079=> "00000000",   --          
-- 0x5A 'Z'        
1080=> "00000000",   --          
1081=> "11111110",   --  ******* 
1082=> "11000110",   --  **   ** 
1083=> "10001100",   --  *   **  
1084=> "00011000",   --     **   
1085=> "00110000",   --    **    
1086=> "01100000",   --   **     
1087=> "11000010",   --  **    * 
1088=> "11000110",   --  **   ** 
1089=> "11111110",   --  ******* 
1090=> "00000000",   --          
1091=> "00000000",   --          
-- 0x5B '['        
1092=> "00000000",   --          
1093=> "01111100",   --   *****  
1094=> "01100000",   --   **     
1095=> "01100000",   --   **     
1096=> "01100000",   --   **     
1097=> "01100000",   --   **     
1098=> "01100000",   --   **     
1099=> "01100000",   --   **     
1100=> "01100000",   --   **     
1101=> "01111100",   --   *****  
1102=> "00000000",   --          
1103=> "00000000",   --          
-- 0x5 C'\'        
1104=> "00000000",   --          
1105=> "00000000",   --          
1106=> "00000000",   --          
1107=> "11000000",   --  **      
1108=> "01100000",   --   **     
1109=> "00110000",   --    **    
1110=> "00011000",   --     **   
1111=> "00001100",   --      **  
1112=> "00000110",   --       ** 
1113=> "00000000",   --          
1114=> "00000000",   --          
1115=> "00000000",   --          
-- 0x5D ']'        
1116=> "00000000",   --          
1117=> "01111100",   --   *****  
1118=> "00001100",   --      **  
1119=> "00001100",   --      **  
1120=> "00001100",   --      **  
1121=> "00001100",   --      **  
1122=> "00001100",   --      **  
1123=> "00001100",   --      **  
1124=> "00001100",   --      **  
1125=> "01111100",   --   *****  
1126=> "00000000",   --          
1127=> "00000000",   --          
-- 0x5E '^'        
1128=> "00000000",   --          
1129=> "00011000",   --     **   
1130=> "00111100",   --    ****  
1131=> "01100110",   --   **  ** 
1132=> "00000000",   --          
1133=> "00000000",   --          
1134=> "00000000",   --          
1135=> "00000000",   --          
1136=> "00000000",   --          
1137=> "00000000",   --          
1138=> "00000000",   --          
1139=> "00000000",   --          
-- 0x5F '_'        
1140=> "00000000",   --          
1141=> "00000000",   --          
1142=> "00000000",   --          
1143=> "00000000",   --          
1144=> "00000000",   --          
1145=> "00000000",   --          
1146=> "00000000",   --          
1147=> "00000000",   --          
1148=> "00000000",   --          
1149=> "00000000",   --          
1150=> "00000000",   --          
1151=> "11111111",   --  ********
-- 0x60 '`'        
1152=> "00011100",   --     ***  
1153=> "00011100",   --     ***  
1154=> "00011000",   --     **   
1155=> "00001100",   --      **  
1156=> "00000000",   --          
1157=> "00000000",   --          
1158=> "00000000",   --          
1159=> "00000000",   --          
1160=> "00000000",   --          
1161=> "00000000",   --          
1162=> "00000000",   --          
1163=> "00000000",   --          
-- 0x61 'a'        
1164=> "00000000",   --          
1165=> "00000000",   --          
1166=> "00000000",   --          
1167=> "00000000",   --          
1168=> "01111000",   --   ****   
1169=> "00001100",   --      **  
1170=> "01111100",   --   *****  
1171=> "11001100",   --  **  **  
1172=> "11011100",   --  ** ***  
1173=> "01110110",   --   *** ** 
1174=> "00000000",   --          
1175=> "00000000",   --          
-- 0x62 'b'        
1176=> "00000000",   --          
1177=> "11100000",   --  ***     
1178=> "01100000",   --   **     
1179=> "01100000",   --   **     
1180=> "01111100",   --   *****  
1181=> "01100110",   --   **  ** 
1182=> "01100110",   --   **  ** 
1183=> "01100110",   --   **  ** 
1184=> "01100110",   --   **  ** 
1185=> "11111100",   --  ******  
1186=> "00000000",   --          
1187=> "00000000",   --          
-- 0x63 'c'        
1188=> "00000000",   --          
1189=> "00000000",   --          
1190=> "00000000",   --          
1191=> "00000000",   --          
1192=> "01111100",   --   *****  
1193=> "11000110",   --  **   ** 
1194=> "11000000",   --  **      
1195=> "11000000",   --  **      
1196=> "11000110",   --  **   ** 
1197=> "01111100",   --   *****  
1198=> "00000000",   --          
1199=> "00000000",   --          
-- 0x64 'd'        
1200=> "00000000",   --          
1201=> "00011100",   --     ***  
1202=> "00001100",   --      **  
1203=> "00001100",   --      **  
1204=> "01111100",   --   *****  
1205=> "11001100",   --  **  **  
1206=> "11001100",   --  **  **  
1207=> "11001100",   --  **  **  
1208=> "11001100",   --  **  **  
1209=> "01111110",   --   ****** 
1210=> "00000000",   --          
1211=> "00000000",   --          
-- 0x65 'e'        
1212=> "00000000",   --          
1213=> "00000000",   --          
1214=> "00000000",   --          
1215=> "00000000",   --          
1216=> "01111100",   --   *****  
1217=> "11000110",   --  **   ** 
1218=> "11111110",   --  ******* 
1219=> "11000000",   --  **      
1220=> "11000110",   --  **   ** 
1221=> "01111100",   --   *****  
1222=> "00000000",   --          
1223=> "00000000",   --          
-- 0x66 'f'        
1224=> "00000000",   --          
1225=> "00011100",   --     ***  
1226=> "00110110",   --    ** ** 
1227=> "00110000",   --    **    
1228=> "00110000",   --    **    
1229=> "11111100",   --  ******  
1230=> "00110000",   --    **    
1231=> "00110000",   --    **    
1232=> "00110000",   --    **    
1233=> "01111000",   --   ****   
1234=> "00000000",   --          
1235=> "00000000",   --          
-- 0x67 'g'        
1236=> "00000000",   --          
1237=> "00000000",   --          
1238=> "00000000",   --          
1239=> "00000000",   --          
1240=> "01110110",   --   *** ** 
1241=> "11001110",   --  **  *** 
1242=> "11000110",   --  **   ** 
1243=> "11000110",   --  **   ** 
1244=> "01111110",   --   ****** 
1245=> "00000110",   --       ** 
1246=> "11000110",   --  **   ** 
1247=> "01111100",   --   *****  
-- 0x68 'h'        
1248=> "00000000",   --          
1249=> "11100000",   --  ***     
1250=> "01100000",   --   **     
1251=> "01100000",   --   **     
1252=> "01101100",   --   ** **  
1253=> "01110110",   --   *** ** 
1254=> "01100110",   --   **  ** 
1255=> "01100110",   --   **  ** 
1256=> "01100110",   --   **  ** 
1257=> "11100110",   --  ***  ** 
1258=> "00000000",   --          
1259=> "00000000",   --          
-- 0x69 'i'        
1260=> "00000000",   --          
1261=> "00011000",   --     **   
1262=> "00011000",   --     **   
1263=> "00000000",   --          
1264=> "00111000",   --    ***   
1265=> "00011000",   --     **   
1266=> "00011000",   --     **   
1267=> "00011000",   --     **   
1268=> "00011000",   --     **   
1269=> "00111100",   --    ****  
1270=> "00000000",   --          
1271=> "00000000",   --          
-- 0x6A 'j'        
1272=> "00000000",   --          
1273=> "00000000",   --          
1274=> "00001100",   --      **  
1275=> "00001100",   --      **  
1276=> "00000000",   --          
1277=> "00011100",   --     ***  
1278=> "00001100",   --      **  
1279=> "00001100",   --      **  
1280=> "00001100",   --      **  
1281=> "11001100",   --  **  **  
1282=> "11001100",   --  **  **  
1283=> "01111000",   --   ****   
-- 0x6B 'k'        
1284=> "00000000",   --          
1285=> "11100000",   --  ***     
1286=> "01100000",   --   **     
1287=> "01100000",   --   **     
1288=> "01100110",   --   **  ** 
1289=> "01101100",   --   ** **  
1290=> "01111000",   --   ****   
1291=> "01101100",   --   ** **  
1292=> "01100110",   --   **  ** 
1293=> "11100110",   --  ***  ** 
1294=> "00000000",   --          
1295=> "00000000",   --          
-- 0x6 C'l'        
1296=> "00000000",   --          
1297=> "01110000",   --   ***    
1298=> "00110000",   --    **    
1299=> "00110000",   --    **    
1300=> "00110000",   --    **    
1301=> "00110000",   --    **    
1302=> "00110000",   --    **    
1303=> "00110000",   --    **    
1304=> "00110100",   --    ** *  
1305=> "00011000",   --     **   
1306=> "00000000",   --          
1307=> "00000000",   --          
-- 0x6D 'm'        
1308=> "00000000",   --          
1309=> "00000000",   --          
1310=> "00000000",   --          
1311=> "00000000",   --          
1312=> "01101100",   --   ** **  
1313=> "11111110",   --  ******* 
1314=> "11010110",   --  ** * ** 
1315=> "11010110",   --  ** * ** 
1316=> "11000110",   --  **   ** 
1317=> "11000110",   --  **   ** 
1318=> "00000000",   --          
1319=> "00000000",   --          
-- 0x6E 'n'        
1320=> "00000000",   --          
1321=> "00000000",   --          
1322=> "00000000",   --          
1323=> "00000000",   --          
1324=> "11011100",   --  ** ***  
1325=> "01100110",   --   **  ** 
1326=> "01100110",   --   **  ** 
1327=> "01100110",   --   **  ** 
1328=> "01100110",   --   **  ** 
1329=> "01100110",   --   **  ** 
1330=> "00000000",   --          
1331=> "00000000",   --          
-- 0x6F 'o'        
1332=> "00000000",   --          
1333=> "00000000",   --          
1334=> "00000000",   --          
1335=> "00000000",   --          
1336=> "01111100",   --   *****  
1337=> "11000110",   --  **   ** 
1338=> "11000110",   --  **   ** 
1339=> "11000110",   --  **   ** 
1340=> "11000110",   --  **   ** 
1341=> "01111100",   --   *****  
1342=> "00000000",   --          
1343=> "00000000",   --          
-- 0x70 'p'        
1344=> "00000000",   --          
1345=> "00000000",   --          
1346=> "00000000",   --          
1347=> "00000000",   --          
1348=> "11011100",   --  ** ***  
1349=> "01100110",   --   **  ** 
1350=> "01100110",   --   **  ** 
1351=> "01100110",   --   **  ** 
1352=> "01111100",   --   *****  
1353=> "01100000",   --   **     
1354=> "01100000",   --   **     
1355=> "11110000",   --  ****    
-- 0x71 'q'        
1356=> "00000000",   --          
1357=> "00000000",   --          
1358=> "00000000",   --          
1359=> "00000000",   --          
1360=> "01110110",   --   *** ** 
1361=> "11001100",   --  **  **  
1362=> "11001100",   --  **  **  
1363=> "11001100",   --  **  **  
1364=> "01111100",   --   *****  
1365=> "00001100",   --      **  
1366=> "00001100",   --      **  
1367=> "00011110",   --     **** 
-- 0x72 'r'        
1368=> "00000000",   --          
1369=> "00000000",   --          
1370=> "00000000",   --          
1371=> "00000000",   --          
1372=> "11011100",   --  ** ***  
1373=> "01100110",   --   **  ** 
1374=> "01100000",   --   **     
1375=> "01100000",   --   **     
1376=> "01100000",   --   **     
1377=> "11110000",   --  ****    
1378=> "00000000",   --          
1379=> "00000000",   --          
-- 0x73 's'        
1380=> "00000000",   --          
1381=> "00000000",   --          
1382=> "00000000",   --          
1383=> "00000000",   --          
1384=> "01111100",   --   *****  
1385=> "11000110",   --  **   ** 
1386=> "01110000",   --   ***    
1387=> "00011100",   --     ***  
1388=> "11000110",   --  **   ** 
1389=> "01111100",   --   *****  
1390=> "00000000",   --          
1391=> "00000000",   --          
-- 0x74 't'        
1392=> "00000000",   --          
1393=> "00110000",   --    **    
1394=> "00110000",   --    **    
1395=> "00110000",   --    **    
1396=> "11111100",   --  ******  
1397=> "00110000",   --    **    
1398=> "00110000",   --    **    
1399=> "00110000",   --    **    
1400=> "00110110",   --    ** ** 
1401=> "00011100",   --     ***  
1402=> "00000000",   --          
1403=> "00000000",   --          
-- 0x75 'u'        
1404=> "00000000",   --          
1405=> "00000000",   --          
1406=> "00000000",   --          
1407=> "00000000",   --          
1408=> "11001100",   --  **  **  
1409=> "11001100",   --  **  **  
1410=> "11001100",   --  **  **  
1411=> "11001100",   --  **  **  
1412=> "11001100",   --  **  **  
1413=> "01110110",   --   *** ** 
1414=> "00000000",   --          
1415=> "00000000",   --          
-- 0x76 'v'        
1416=> "00000000",   --          
1417=> "00000000",   --          
1418=> "00000000",   --          
1419=> "00000000",   --          
1420=> "11000110",   --  **   ** 
1421=> "11000110",   --  **   ** 
1422=> "11000110",   --  **   ** 
1423=> "01101100",   --   ** **  
1424=> "00111000",   --    ***   
1425=> "00010000",   --     *    
1426=> "00000000",   --          
1427=> "00000000",   --          
-- 0x77 'w'        
1428=> "00000000",   --          
1429=> "00000000",   --          
1430=> "00000000",   --          
1431=> "00000000",   --          
1432=> "11000110",   --  **   ** 
1433=> "11000110",   --  **   ** 
1434=> "11010110",   --  ** * ** 
1435=> "11010110",   --  ** * ** 
1436=> "11111110",   --  ******* 
1437=> "01101100",   --   ** **  
1438=> "00000000",   --          
1439=> "00000000",   --          
-- 0x78 'x'        
1440=> "00000000",   --          
1441=> "00000000",   --          
1442=> "00000000",   --          
1443=> "00000000",   --          
1444=> "11000110",   --  **   ** 
1445=> "01101100",   --   ** **  
1446=> "00111000",   --    ***   
1447=> "00111000",   --    ***   
1448=> "01101100",   --   ** **  
1449=> "11000110",   --  **   ** 
1450=> "00000000",   --          
1451=> "00000000",   --          
-- 0x79 'y'        
1452=> "00000000",   --          
1453=> "00000000",   --          
1454=> "00000000",   --          
1455=> "00000000",   --          
1456=> "11000110",   --  **   ** 
1457=> "11000110",   --  **   ** 
1458=> "11000110",   --  **   ** 
1459=> "11001110",   --  **  *** 
1460=> "01110110",   --   *** ** 
1461=> "00000110",   --       ** 
1462=> "11000110",   --  **   ** 
1463=> "01111100",   --   *****  
-- 0x7A 'z'        
1464=> "00000000",   --          
1465=> "00000000",   --          
1466=> "00000000",   --          
1467=> "00000000",   --          
1468=> "11111110",   --  ******* 
1469=> "10001100",   --  *   **  
1470=> "00011000",   --     **   
1471=> "00110000",   --    **    
1472=> "01100010",   --   **   * 
1473=> "11111110",   --  ******* 
1474=> "00000000",   --          
1475=> "00000000",   --          
-- 0x7B '{'        
1476=> "00000000",   --          
1477=> "00001110",   --      *** 
1478=> "00011000",   --     **   
1479=> "00011000",   --     **   
1480=> "00011000",   --     **   
1481=> "01110000",   --   ***    
1482=> "00011000",   --     **   
1483=> "00011000",   --     **   
1484=> "00011000",   --     **   
1485=> "00001110",   --      *** 
1486=> "00000000",   --          
1487=> "00000000",   --          
-- 0x7 C'|'        
1488=> "00000000",   --          
1489=> "00011000",   --     **   
1490=> "00011000",   --     **   
1491=> "00011000",   --     **   
1492=> "00011000",   --     **   
1493=> "00011000",   --     **   
1494=> "00011000",   --     **   
1495=> "00011000",   --     **   
1496=> "00011000",   --     **   
1497=> "00011000",   --     **   
1498=> "00000000",   --          
1499=> "00000000",   --          
-- 0x7D '}'        
1500=> "00000000",   --          
1501=> "01110000",   --   ***    
1502=> "00011000",   --     **   
1503=> "00011000",   --     **   
1504=> "00011000",   --     **   
1505=> "00001110",   --      *** 
1506=> "00011000",   --     **   
1507=> "00011000",   --     **   
1508=> "00011000",   --     **   
1509=> "01110000",   --   ***    
1510=> "00000000",   --          
1511=> "00000000",   --          
-- 0x7E '~'        
1512=> "00000000",   --          
1513=> "01110110",   --   *** ** 
1514=> "11011100",   --  ** ***  
1515=> "00000000",   --          
1516=> "00000000",   --          
1517=> "00000000",   --          
1518=> "00000000",   --          
1519=> "00000000",   --          
1520=> "00000000",   --          
1521=> "00000000",   --          
1522=> "00000000",   --          
1523=> "00000000",   --          
-- 0x7F ''         
1524=> "01100110",   --   **  ** 
1525=> "01100110",   --   **  ** 
1526=> "00000000",   --          
1527=> "01100110",   --   **  ** 
1528=> "01100110",   --   **  ** 
1529=> "01100110",   --   **  ** 
1530=> "00111100",   --    ****  
1531=> "00011000",   --     **   
1532=> "00011000",   --     **   
1533=> "00111100",   --    ****  
1534=> "00000000",   --          
1535=> "00000000",   --          
-- 0x80 ''         
1536=> "00110000",   --    **    
1537=> "00011000",   --     **   
1538=> "00000000",   --          
1539=> "00111000",   --    ***   
1540=> "01101100",   --   ** **  
1541=> "11000110",   --  **   ** 
1542=> "11000110",   --  **   ** 
1543=> "11111110",   --  ******* 
1544=> "11000110",   --  **   ** 
1545=> "11000110",   --  **   ** 
1546=> "00000000",   --          
1547=> "00000000",   --          
-- 0x81 ''         
1548=> "00011000",   --     **   
1549=> "00110000",   --    **    
1550=> "00000000",   --          
1551=> "00111000",   --    ***   
1552=> "01101100",   --   ** **  
1553=> "11000110",   --  **   ** 
1554=> "11000110",   --  **   ** 
1555=> "11111110",   --  ******* 
1556=> "11000110",   --  **   ** 
1557=> "11000110",   --  **   ** 
1558=> "00000000",   --          
1559=> "00000000",   --          
-- 0x82 ''         
1560=> "00111000",   --    ***   
1561=> "01101100",   --   ** **  
1562=> "00111000",   --    ***   
1563=> "00000000",   --          
1564=> "01111100",   --   *****  
1565=> "11000110",   --  **   ** 
1566=> "11000110",   --  **   ** 
1567=> "11111110",   --  ******* 
1568=> "11000110",   --  **   ** 
1569=> "11000110",   --  **   ** 
1570=> "00000000",   --          
1571=> "00000000",   --          
-- 0x83 ''         
1572=> "01110110",   --   *** ** 
1573=> "11011100",   --  ** ***  
1574=> "00000000",   --          
1575=> "00111000",   --    ***   
1576=> "01101100",   --   ** **  
1577=> "11000110",   --  **   ** 
1578=> "11000110",   --  **   ** 
1579=> "11111110",   --  ******* 
1580=> "11000110",   --  **   ** 
1581=> "11000110",   --  **   ** 
1582=> "00000000",   --          
1583=> "00000000",   --          
-- 0x84 ''         
1584=> "01101100",   --   ** **  
1585=> "01101100",   --   ** **  
1586=> "00000000",   --          
1587=> "00111000",   --    ***   
1588=> "01101100",   --   ** **  
1589=> "11000110",   --  **   ** 
1590=> "11000110",   --  **   ** 
1591=> "11111110",   --  ******* 
1592=> "11000110",   --  **   ** 
1593=> "11000110",   --  **   ** 
1594=> "00000000",   --          
1595=> "00000000",   --          
-- 0x85 ''         
1596=> "00111000",   --    ***   
1597=> "01101100",   --   ** **  
1598=> "00111000",   --    ***   
1599=> "00000000",   --          
1600=> "01111100",   --   *****  
1601=> "11000110",   --  **   ** 
1602=> "11000110",   --  **   ** 
1603=> "11111110",   --  ******* 
1604=> "11000110",   --  **   ** 
1605=> "11000110",   --  **   ** 
1606=> "00000000",   --          
1607=> "00000000",   --          
-- 0x86 ''         
1608=> "01111110",   --   ****** 
1609=> "11011000",   --  ** **   
1610=> "11011000",   --  ** **   
1611=> "11011000",   --  ** **   
1612=> "11011000",   --  ** **   
1613=> "11111110",   --  ******* 
1614=> "11011000",   --  ** **   
1615=> "11011000",   --  ** **   
1616=> "11011000",   --  ** **   
1617=> "11011110",   --  ** **** 
1618=> "00000000",   --          
1619=> "00000000",   --          
-- 0x87 ''         
1620=> "00000000",   --          
1621=> "00111100",   --    ****  
1622=> "01100110",   --   **  ** 
1623=> "11000000",   --  **      
1624=> "11000000",   --  **      
1625=> "11000000",   --  **      
1626=> "11000110",   --  **   ** 
1627=> "01100110",   --   **  ** 
1628=> "00111100",   --    ****  
1629=> "00011000",   --     **   
1630=> "11001100",   --  **  **  
1631=> "00111000",   --    ***   
-- 0x88 ''         
1632=> "00011000",   --     **   
1633=> "00001100",   --      **  
1634=> "00000000",   --          
1635=> "11111110",   --  ******* 
1636=> "01100110",   --   **  ** 
1637=> "01100000",   --   **     
1638=> "01111100",   --   *****  
1639=> "01100000",   --   **     
1640=> "01100110",   --   **  ** 
1641=> "11111110",   --  ******* 
1642=> "00000000",   --          
1643=> "00000000",   --          
-- 0x89 ''         
1644=> "00011000",   --     **   
1645=> "00110000",   --    **    
1646=> "00000000",   --          
1647=> "11111110",   --  ******* 
1648=> "01100110",   --   **  ** 
1649=> "01100000",   --   **     
1650=> "01111100",   --   *****  
1651=> "01100000",   --   **     
1652=> "01100110",   --   **  ** 
1653=> "11111110",   --  ******* 
1654=> "00000000",   --          
1655=> "00000000",   --          
-- 0x8A ''         
1656=> "00111000",   --    ***   
1657=> "01101100",   --   ** **  
1658=> "00000000",   --          
1659=> "11111110",   --  ******* 
1660=> "01100110",   --   **  ** 
1661=> "01100000",   --   **     
1662=> "01111100",   --   *****  
1663=> "01100000",   --   **     
1664=> "01100110",   --   **  ** 
1665=> "11111110",   --  ******* 
1666=> "00000000",   --          
1667=> "00000000",   --          
-- 0x8B ''         
1668=> "01101100",   --   ** **  
1669=> "01101100",   --   ** **  
1670=> "00000000",   --          
1671=> "11111110",   --  ******* 
1672=> "01100110",   --   **  ** 
1673=> "01100000",   --   **     
1674=> "01111100",   --   *****  
1675=> "01100000",   --   **     
1676=> "01100110",   --   **  ** 
1677=> "11111110",   --  ******* 
1678=> "00000000",   --          
1679=> "00000000",   --          
-- 0x8 C''         
1680=> "00011000",   --     **   
1681=> "00001100",   --      **  
1682=> "00000000",   --          
1683=> "00111100",   --    ****  
1684=> "00011000",   --     **   
1685=> "00011000",   --     **   
1686=> "00011000",   --     **   
1687=> "00011000",   --     **   
1688=> "00011000",   --     **   
1689=> "00111100",   --    ****  
1690=> "00000000",   --          
1691=> "00000000",   --          
-- 0x8D ''         
1692=> "00011000",   --     **   
1693=> "00110000",   --    **    
1694=> "00000000",   --          
1695=> "00111100",   --    ****  
1696=> "00011000",   --     **   
1697=> "00011000",   --     **   
1698=> "00011000",   --     **   
1699=> "00011000",   --     **   
1700=> "00011000",   --     **   
1701=> "00111100",   --    ****  
1702=> "00000000",   --          
1703=> "00000000",   --          
-- 0x8E ''         
1704=> "00111100",   --    ****  
1705=> "01100110",   --   **  ** 
1706=> "00000000",   --          
1707=> "00111100",   --    ****  
1708=> "00011000",   --     **   
1709=> "00011000",   --     **   
1710=> "00011000",   --     **   
1711=> "00011000",   --     **   
1712=> "00011000",   --     **   
1713=> "00111100",   --    ****  
1714=> "00000000",   --          
1715=> "00000000",   --          
-- 0x8F ''         
1716=> "01100110",   --   **  ** 
1717=> "01100110",   --   **  ** 
1718=> "00000000",   --          
1719=> "00111100",   --    ****  
1720=> "00011000",   --     **   
1721=> "00011000",   --     **   
1722=> "00011000",   --     **   
1723=> "00011000",   --     **   
1724=> "00011000",   --     **   
1725=> "00111100",   --    ****  
1726=> "00000000",   --          
1727=> "00000000",   --          
-- 0x90 ''         
1728=> "00000000",   --          
1729=> "11111000",   --  *****   
1730=> "01101100",   --   ** **  
1731=> "01100110",   --   **  ** 
1732=> "01100110",   --   **  ** 
1733=> "11110110",   --  **** ** 
1734=> "01100110",   --   **  ** 
1735=> "01100110",   --   **  ** 
1736=> "01101100",   --   ** **  
1737=> "11111000",   --  *****   
1738=> "00000000",   --          
1739=> "00000000",   --          
-- 0x91 ''         
1740=> "01110110",   --   *** ** 
1741=> "11011100",   --  ** ***  
1742=> "00000000",   --          
1743=> "11000110",   --  **   ** 
1744=> "11100110",   --  ***  ** 
1745=> "11110110",   --  **** ** 
1746=> "11011110",   --  ** **** 
1747=> "11001110",   --  **  *** 
1748=> "11000110",   --  **   ** 
1749=> "11000110",   --  **   ** 
1750=> "00000000",   --          
1751=> "00000000",   --          
-- 0x92 ''         
1752=> "00110000",   --    **    
1753=> "00011000",   --     **   
1754=> "00000000",   --          
1755=> "01111100",   --   *****  
1756=> "11000110",   --  **   ** 
1757=> "11000110",   --  **   ** 
1758=> "11000110",   --  **   ** 
1759=> "11000110",   --  **   ** 
1760=> "11000110",   --  **   ** 
1761=> "01111100",   --   *****  
1762=> "00000000",   --          
1763=> "00000000",   --          
-- 0x93 ''         
1764=> "00011000",   --     **   
1765=> "00110000",   --    **    
1766=> "00000000",   --          
1767=> "01111100",   --   *****  
1768=> "11000110",   --  **   ** 
1769=> "11000110",   --  **   ** 
1770=> "11000110",   --  **   ** 
1771=> "11000110",   --  **   ** 
1772=> "11000110",   --  **   ** 
1773=> "01111100",   --   *****  
1774=> "00000000",   --          
1775=> "00000000",   --          
-- 0x94 ''         
1776=> "00111000",   --    ***   
1777=> "01101100",   --   ** **  
1778=> "00000000",   --          
1779=> "01111100",   --   *****  
1780=> "11000110",   --  **   ** 
1781=> "11000110",   --  **   ** 
1782=> "11000110",   --  **   ** 
1783=> "11000110",   --  **   ** 
1784=> "11000110",   --  **   ** 
1785=> "01111100",   --   *****  
1786=> "00000000",   --          
1787=> "00000000",   --          
-- 0x95 ''         
1788=> "01110110",   --   *** ** 
1789=> "11011100",   --  ** ***  
1790=> "00000000",   --          
1791=> "01111100",   --   *****  
1792=> "11000110",   --  **   ** 
1793=> "11000110",   --  **   ** 
1794=> "11000110",   --  **   ** 
1795=> "11000110",   --  **   ** 
1796=> "11000110",   --  **   ** 
1797=> "01111100",   --   *****  
1798=> "00000000",   --          
1799=> "00000000",   --          
-- 0x96 ''         
1800=> "01101100",   --   ** **  
1801=> "01101100",   --   ** **  
1802=> "00000000",   --          
1803=> "01111100",   --   *****  
1804=> "11000110",   --  **   ** 
1805=> "11000110",   --  **   ** 
1806=> "11000110",   --  **   ** 
1807=> "11000110",   --  **   ** 
1808=> "11000110",   --  **   ** 
1809=> "01111100",   --   *****  
1810=> "00000000",   --          
1811=> "00000000",   --          
-- 0x97 ''         
1812=> "00000000",   --          
1813=> "00000000",   --          
1814=> "00000000",   --          
1815=> "00000000",   --          
1816=> "01101100",   --   ** **  
1817=> "00111000",   --    ***   
1818=> "00111000",   --    ***   
1819=> "01101100",   --   ** **  
1820=> "00000000",   --          
1821=> "00000000",   --          
1822=> "00000000",   --          
1823=> "00000000",   --          
-- 0x98 ''         
1824=> "00000000",   --          
1825=> "01111110",   --   ****** 
1826=> "11000110",   --  **   ** 
1827=> "11001110",   --  **  *** 
1828=> "11011110",   --  ** **** 
1829=> "11010110",   --  ** * ** 
1830=> "11110110",   --  **** ** 
1831=> "11100110",   --  ***  ** 
1832=> "11000110",   --  **   ** 
1833=> "11111100",   --  ******  
1834=> "00000000",   --          
1835=> "00000000",   --          
-- 0x99 ''         
1836=> "00110000",   --    **    
1837=> "00011000",   --     **   
1838=> "00000000",   --          
1839=> "11000110",   --  **   ** 
1840=> "11000110",   --  **   ** 
1841=> "11000110",   --  **   ** 
1842=> "11000110",   --  **   ** 
1843=> "11000110",   --  **   ** 
1844=> "11000110",   --  **   ** 
1845=> "01111100",   --   *****  
1846=> "00000000",   --          
1847=> "00000000",   --          
-- 0x9A ''         
1848=> "00011000",   --     **   
1849=> "00110000",   --    **    
1850=> "00000000",   --          
1851=> "11000110",   --  **   ** 
1852=> "11000110",   --  **   ** 
1853=> "11000110",   --  **   ** 
1854=> "11000110",   --  **   ** 
1855=> "11000110",   --  **   ** 
1856=> "11000110",   --  **   ** 
1857=> "01111100",   --   *****  
1858=> "00000000",   --          
1859=> "00000000",   --          
-- 0x9B ''         
1860=> "00111000",   --    ***   
1861=> "01101100",   --   ** **  
1862=> "00000000",   --          
1863=> "11000110",   --  **   ** 
1864=> "11000110",   --  **   ** 
1865=> "11000110",   --  **   ** 
1866=> "11000110",   --  **   ** 
1867=> "11000110",   --  **   ** 
1868=> "11000110",   --  **   ** 
1869=> "01111100",   --   *****  
1870=> "00000000",   --          
1871=> "00000000",   --          
-- 0x9 C''         
1872=> "01101100",   --   ** **  
1873=> "01101100",   --   ** **  
1874=> "00000000",   --          
1875=> "11000110",   --  **   ** 
1876=> "11000110",   --  **   ** 
1877=> "11000110",   --  **   ** 
1878=> "11000110",   --  **   ** 
1879=> "11000110",   --  **   ** 
1880=> "11000110",   --  **   ** 
1881=> "01111100",   --   *****  
1882=> "00000000",   --          
1883=> "00000000",   --          
-- 0x9D ''         
1884=> "00001100",   --      **  
1885=> "00011000",   --     **   
1886=> "00000000",   --          
1887=> "01100110",   --   **  ** 
1888=> "01100110",   --   **  ** 
1889=> "01100110",   --   **  ** 
1890=> "00111100",   --    ****  
1891=> "00011000",   --     **   
1892=> "00011000",   --     **   
1893=> "00111100",   --    ****  
1894=> "00000000",   --          
1895=> "00000000",   --          
-- 0x9E ''         
1896=> "00000000",   --          
1897=> "11110000",   --  ****    
1898=> "01100000",   --   **     
1899=> "01111100",   --   *****  
1900=> "01100110",   --   **  ** 
1901=> "01100110",   --   **  ** 
1902=> "01100110",   --   **  ** 
1903=> "01111100",   --   *****  
1904=> "01100000",   --   **     
1905=> "11110000",   --  ****    
1906=> "00000000",   --          
1907=> "00000000",   --          
-- 0x9F ''         
1908=> "00000000",   --          
1909=> "01111100",   --   *****  
1910=> "11000110",   --  **   ** 
1911=> "11000110",   --  **   ** 
1912=> "11000110",   --  **   ** 
1913=> "11001100",   --  **  **  
1914=> "11000110",   --  **   ** 
1915=> "11000110",   --  **   ** 
1916=> "11010110",   --  ** * ** 
1917=> "11011100",   --  ** ***  
1918=> "10000000",   --  *       
1919=> "00000000",   --          
-- 0xA0 ''         
1920=> "00000000",   --          
1921=> "00000000",   --          
1922=> "00000000",   --          
1923=> "00000000",   --          
1924=> "00000000",   --          
1925=> "00000000",   --          
1926=> "00000000",   --          
1927=> "00000000",   --          
1928=> "00000000",   --          
1929=> "10000010",   --  *     * 
1930=> "11111110",   --  ******* 
1931=> "00000000",   --          
-- 0xA1 ''         
1932=> "00000000",   --          
1933=> "00000000",   --          
1934=> "00000000",   --          
1935=> "00011000",   --     **   
1936=> "00011000",   --     **   
1937=> "00000000",   --          
1938=> "00011000",   --     **   
1939=> "00011000",   --     **   
1940=> "00111100",   --    ****  
1941=> "00111100",   --    ****  
1942=> "00111100",   --    ****  
1943=> "00011000",   --     **   
-- 0xA2 ''         
1944=> "00000000",   --          
1945=> "00000000",   --          
1946=> "00010000",   --     *    
1947=> "01111100",   --   *****  
1948=> "11010110",   --  ** * ** 
1949=> "11010000",   --  ** *    
1950=> "11010000",   --  ** *    
1951=> "11010110",   --  ** * ** 
1952=> "01111100",   --   *****  
1953=> "00010000",   --     *    
1954=> "00000000",   --          
1955=> "00000000",   --          
-- 0xA3 ''         
1956=> "00000000",   --          
1957=> "00111000",   --    ***   
1958=> "01101100",   --   ** **  
1959=> "01100000",   --   **     
1960=> "01100000",   --   **     
1961=> "11110000",   --  ****    
1962=> "01100000",   --   **     
1963=> "01100110",   --   **  ** 
1964=> "11110110",   --  **** ** 
1965=> "01101100",   --   ** **  
1966=> "00000000",   --          
1967=> "00000000",   --          
-- 0xA4 ''         
1968=> "00000000",   --          
1969=> "00111100",   --    ****  
1970=> "01100010",   --   **   * 
1971=> "01100000",   --   **     
1972=> "11111000",   --  *****   
1973=> "01100000",   --   **     
1974=> "11111000",   --  *****   
1975=> "01100000",   --   **     
1976=> "01100010",   --   **   * 
1977=> "00111100",   --    ****  
1978=> "00000000",   --          
1979=> "00000000",   --          
-- 0xA5 ''         
1980=> "00000000",   --          
1981=> "01100110",   --   **  ** 
1982=> "01100110",   --   **  ** 
1983=> "00111100",   --    ****  
1984=> "00011000",   --     **   
1985=> "01111110",   --   ****** 
1986=> "00011000",   --     **   
1987=> "00111100",   --    ****  
1988=> "00011000",   --     **   
1989=> "00011000",   --     **   
1990=> "00000000",   --          
1991=> "00000000",   --          
-- 0xA6 ''         
1992=> "01101100",   --   ** **  
1993=> "00111000",   --    ***   
1994=> "00000000",   --          
1995=> "01111100",   --   *****  
1996=> "11000110",   --  **   ** 
1997=> "11000000",   --  **      
1998=> "01111100",   --   *****  
1999=> "00000110",   --       ** 
2000=> "11000110",   --  **   ** 
2001=> "01111100",   --   *****  
2002=> "00000000",   --          
2003=> "00000000",   --          
-- 0xA7 ''         
2004=> "01111100",   --   *****  
2005=> "11000110",   --  **   ** 
2006=> "11000110",   --  **   ** 
2007=> "01100000",   --   **     
2008=> "01111100",   --   *****  
2009=> "11000110",   --  **   ** 
2010=> "11000110",   --  **   ** 
2011=> "01111100",   --   *****  
2012=> "00001100",   --      **  
2013=> "11000110",   --  **   ** 
2014=> "11000110",   --  **   ** 
2015=> "01111100",   --   *****  
-- 0xA8 ''         
2016=> "00000000",   --          
2017=> "01101100",   --   ** **  
2018=> "00111000",   --    ***   
2019=> "00000000",   --          
2020=> "01111100",   --   *****  
2021=> "11000110",   --  **   ** 
2022=> "01110000",   --   ***    
2023=> "00011100",   --     ***  
2024=> "11000110",   --  **   ** 
2025=> "01111100",   --   *****  
2026=> "00000000",   --          
2027=> "00000000",   --          
-- 0xA9 ''         
2028=> "01111110",   --   ****** 
2029=> "10000001",   --  *      *
2030=> "10011001",   --  *  **  *
2031=> "10100101",   --  * *  * *
2032=> "10100001",   --  * *    *
2033=> "10100001",   --  * *    *
2034=> "10100101",   --  * *  * *
2035=> "10011001",   --  *  **  *
2036=> "10000001",   --  *      *
2037=> "01111110",   --   ****** 
2038=> "00000000",   --          
2039=> "00000000",   --          
-- 0xAA ''         
2040=> "00111100",   --    ****  
2041=> "01101100",   --   ** **  
2042=> "01101100",   --   ** **  
2043=> "00111110",   --    ***** 
2044=> "00000000",   --          
2045=> "01111110",   --   ****** 
2046=> "00000000",   --          
2047=> "00000000",   --          
2048=> "00000000",   --          
2049=> "00000000",   --          
2050=> "00000000",   --          
2051=> "00000000",   --          
-- 0xAB ''         
2052=> "00000000",   --          
2053=> "00000000",   --          
2054=> "00000000",   --          
2055=> "00110110",   --    ** ** 
2056=> "01101100",   --   ** **  
2057=> "11011000",   --  ** **   
2058=> "01101100",   --   ** **  
2059=> "00110110",   --    ** ** 
2060=> "00000000",   --          
2061=> "00000000",   --          
2062=> "00000000",   --          
2063=> "00000000",   --          
-- 0xA C''         
2064=> "00000000",   --          
2065=> "00000000",   --          
2066=> "00000000",   --          
2067=> "00000000",   --          
2068=> "00000000",   --          
2069=> "01111110",   --   ****** 
2070=> "00000110",   --       ** 
2071=> "00000110",   --       ** 
2072=> "00000110",   --       ** 
2073=> "00000000",   --          
2074=> "00000000",   --          
2075=> "00000000",   --          
-- 0xAD ''         
2076=> "00000000",   --          
2077=> "00000000",   --          
2078=> "00000000",   --          
2079=> "00000000",   --          
2080=> "00000000",   --          
2081=> "01111110",   --   ****** 
2082=> "00000000",   --          
2083=> "00000000",   --          
2084=> "00000000",   --          
2085=> "00000000",   --          
2086=> "00000000",   --          
2087=> "00000000",   --          
-- 0xAE ''         
2088=> "01111110",   --   ****** 
2089=> "10000001",   --  *      *
2090=> "10111001",   --  * ***  *
2091=> "10100101",   --  * *  * *
2092=> "10100101",   --  * *  * *
2093=> "10111001",   --  * ***  *
2094=> "10100101",   --  * *  * *
2095=> "10100101",   --  * *  * *
2096=> "10000001",   --  *      *
2097=> "01111110",   --   ****** 
2098=> "00000000",   --          
2099=> "00000000",   --          
-- 0xAF ''         
2100=> "11111111",   --  ********
2101=> "00000000",   --          
2102=> "00000000",   --          
2103=> "00000000",   --          
2104=> "00000000",   --          
2105=> "00000000",   --          
2106=> "00000000",   --          
2107=> "00000000",   --          
2108=> "00000000",   --          
2109=> "00000000",   --          
2110=> "00000000",   --          
2111=> "00000000",   --          
-- 0xB0 ''         
2112=> "00000000",   --          
2113=> "00111000",   --    ***   
2114=> "01101100",   --   ** **  
2115=> "00111000",   --    ***   
2116=> "00000000",   --          
2117=> "00000000",   --          
2118=> "00000000",   --          
2119=> "00000000",   --          
2120=> "00000000",   --          
2121=> "00000000",   --          
2122=> "00000000",   --          
2123=> "00000000",   --          
-- 0xB1 ''         
2124=> "00000000",   --          
2125=> "00000000",   --          
2126=> "00000000",   --          
2127=> "00011000",   --     **   
2128=> "00011000",   --     **   
2129=> "01111110",   --   ****** 
2130=> "00011000",   --     **   
2131=> "00011000",   --     **   
2132=> "00000000",   --          
2133=> "01111110",   --   ****** 
2134=> "00000000",   --          
2135=> "00000000",   --          
-- 0xB2 ''         
2136=> "00000000",   --          
2137=> "00111000",   --    ***   
2138=> "01101100",   --   ** **  
2139=> "00011000",   --     **   
2140=> "00110000",   --    **    
2141=> "01111100",   --   *****  
2142=> "00000000",   --          
2143=> "00000000",   --          
2144=> "00000000",   --          
2145=> "00000000",   --          
2146=> "00000000",   --          
2147=> "00000000",   --          
-- 0xB3 ''         
2148=> "00000000",   --          
2149=> "00111000",   --    ***   
2150=> "01101100",   --   ** **  
2151=> "00011000",   --     **   
2152=> "01101100",   --   ** **  
2153=> "00111000",   --    ***   
2154=> "00000000",   --          
2155=> "00000000",   --          
2156=> "00000000",   --          
2157=> "00000000",   --          
2158=> "00000000",   --          
2159=> "00000000",   --          
-- 0xB4 ''         
2160=> "01101100",   --   ** **  
2161=> "00111000",   --    ***   
2162=> "00000000",   --          
2163=> "11111110",   --  ******* 
2164=> "11000110",   --  **   ** 
2165=> "00001100",   --      **  
2166=> "00111000",   --    ***   
2167=> "01100010",   --   **   * 
2168=> "11000110",   --  **   ** 
2169=> "11111110",   --  ******* 
2170=> "00000000",   --          
2171=> "00000000",   --          
-- 0xB5 ''         
2172=> "00000000",   --          
2173=> "00000000",   --          
2174=> "00000000",   --          
2175=> "00000000",   --          
2176=> "11001100",   --  **  **  
2177=> "11001100",   --  **  **  
2178=> "11001100",   --  **  **  
2179=> "11001100",   --  **  **  
2180=> "11001100",   --  **  **  
2181=> "11110110",   --  **** ** 
2182=> "11000000",   --  **      
2183=> "11000000",   --  **      
-- 0xB6 ''         
2184=> "00000000",   --          
2185=> "01111111",   --   *******
2186=> "11011011",   --  ** ** **
2187=> "11011011",   --  ** ** **
2188=> "11011011",   --  ** ** **
2189=> "01111011",   --   **** **
2190=> "00011011",   --     ** **
2191=> "00011011",   --     ** **
2192=> "00011011",   --     ** **
2193=> "00011011",   --     ** **
2194=> "00000000",   --          
2195=> "00000000",   --          
-- 0xB7 ''         
2196=> "00000000",   --          
2197=> "00000000",   --          
2198=> "00000000",   --          
2199=> "00000000",   --          
2200=> "00000000",   --          
2201=> "00011000",   --     **   
2202=> "00011000",   --     **   
2203=> "00000000",   --          
2204=> "00000000",   --          
2205=> "00000000",   --          
2206=> "00000000",   --          
2207=> "00000000",   --          
-- 0xB8 ''         
2208=> "00000000",   --          
2209=> "01101100",   --   ** **  
2210=> "00111000",   --    ***   
2211=> "00000000",   --          
2212=> "11111110",   --  ******* 
2213=> "10001100",   --  *   **  
2214=> "00011000",   --     **   
2215=> "00110000",   --    **    
2216=> "01100010",   --   **   * 
2217=> "11111110",   --  ******* 
2218=> "00000000",   --          
2219=> "00000000",   --          
-- 0xB9 ''         
2220=> "00000000",   --          
2221=> "00110000",   --    **    
2222=> "01110000",   --   ***    
2223=> "00110000",   --    **    
2224=> "00110000",   --    **    
2225=> "01111000",   --   ****   
2226=> "00000000",   --          
2227=> "00000000",   --          
2228=> "00000000",   --          
2229=> "00000000",   --          
2230=> "00000000",   --          
2231=> "00000000",   --          
-- 0xBA ''         
2232=> "00111000",   --    ***   
2233=> "01101100",   --   ** **  
2234=> "01101100",   --   ** **  
2235=> "00111000",   --    ***   
2236=> "00000000",   --          
2237=> "01111100",   --   *****  
2238=> "00000000",   --          
2239=> "00000000",   --          
2240=> "00000000",   --          
2241=> "00000000",   --          
2242=> "00000000",   --          
2243=> "00000000",   --          
-- 0xBB ''         
2244=> "00000000",   --          
2245=> "00000000",   --          
2246=> "00000000",   --          
2247=> "11011000",   --  ** **   
2248=> "01101100",   --   ** **  
2249=> "00110110",   --    ** ** 
2250=> "01101100",   --   ** **  
2251=> "11011000",   --  ** **   
2252=> "00000000",   --          
2253=> "00000000",   --          
2254=> "00000000",   --          
2255=> "00000000",   --          
-- 0xB C''         
2256=> "00000000",   --          
2257=> "01101110",   --   ** *** 
2258=> "11011011",   --  ** ** **
2259=> "11011011",   --  ** ** **
2260=> "11011111",   --  ** *****
2261=> "11011000",   --  ** **   
2262=> "11011000",   --  ** **   
2263=> "11011001",   --  ** **  *
2264=> "11011111",   --  ** *****
2265=> "01101110",   --   ** *** 
2266=> "00000000",   --          
2267=> "00000000",   --          
-- 0xBD ''         
2268=> "00000000",   --          
2269=> "00000000",   --          
2270=> "00000000",   --          
2271=> "00000000",   --          
2272=> "01101100",   --   ** **  
2273=> "11011010",   --  ** ** * 
2274=> "11011110",   --  ** **** 
2275=> "11011000",   --  ** **   
2276=> "11011010",   --  ** ** * 
2277=> "01101100",   --   ** **  
2278=> "00000000",   --          
2279=> "00000000",   --          
-- 0xBE ''         
2280=> "01100110",   --   **  ** 
2281=> "01100110",   --   **  ** 
2282=> "00000000",   --          
2283=> "01100110",   --   **  ** 
2284=> "01100110",   --   **  ** 
2285=> "00111100",   --    ****  
2286=> "00011000",   --     **   
2287=> "00011000",   --     **   
2288=> "00011000",   --     **   
2289=> "00111100",   --    ****  
2290=> "00000000",   --          
2291=> "00000000",   --          
-- 0xBF ''         
2292=> "00000000",   --          
2293=> "00000000",   --          
2294=> "00000000",   --          
2295=> "00110000",   --    **    
2296=> "00110000",   --    **    
2297=> "00000000",   --          
2298=> "00110000",   --    **    
2299=> "00110000",   --    **    
2300=> "01100000",   --   **     
2301=> "11000110",   --  **   ** 
2302=> "11000110",   --  **   ** 
2303=> "01111100",   --   *****  
-- 0xC0 ''         
2304=> "00000000",   --          
2305=> "00000000",   --          
2306=> "11111111",   --  ********
2307=> "00000000",   --          
2308=> "00000000",   --          
2309=> "00000000",   --          
2310=> "00000000",   --          
2311=> "00000000",   --          
2312=> "00000000",   --          
2313=> "00000000",   --          
2314=> "00000000",   --          
2315=> "00000000",   --          
-- 0xC1 ''         
2316=> "00011000",   --     **   
2317=> "00011000",   --     **   
2318=> "00011000",   --     **   
2319=> "00011000",   --     **   
2320=> "00011000",   --     **   
2321=> "00011000",   --     **   
2322=> "00000000",   --          
2323=> "00000000",   --          
2324=> "00000000",   --          
2325=> "00000000",   --          
2326=> "00000000",   --          
2327=> "00000000",   --          
-- 0xC2 ''         
2328=> "00000000",   --          
2329=> "00000000",   --          
2330=> "00000000",   --          
2331=> "00000000",   --          
2332=> "00000000",   --          
2333=> "00011111",   --     *****
2334=> "00000000",   --          
2335=> "00000000",   --          
2336=> "00000000",   --          
2337=> "00000000",   --          
2338=> "00000000",   --          
2339=> "00000000",   --          
-- 0xC3 ''         
2340=> "00011000",   --     **   
2341=> "00011000",   --     **   
2342=> "00011000",   --     **   
2343=> "00011000",   --     **   
2344=> "00011000",   --     **   
2345=> "00011111",   --     *****
2346=> "00000000",   --          
2347=> "00000000",   --          
2348=> "00000000",   --          
2349=> "00000000",   --          
2350=> "00000000",   --          
2351=> "00000000",   --          
-- 0xC4 ''         
2352=> "00000000",   --          
2353=> "00000000",   --          
2354=> "00000000",   --          
2355=> "00000000",   --          
2356=> "00000000",   --          
2357=> "00011000",   --     **   
2358=> "00011000",   --     **   
2359=> "00011000",   --     **   
2360=> "00011000",   --     **   
2361=> "00011000",   --     **   
2362=> "00011000",   --     **   
2363=> "00011000",   --     **   
-- 0xC5 ''         
2364=> "00011000",   --     **   
2365=> "00011000",   --     **   
2366=> "00011000",   --     **   
2367=> "00011000",   --     **   
2368=> "00011000",   --     **   
2369=> "00011000",   --     **   
2370=> "00011000",   --     **   
2371=> "00011000",   --     **   
2372=> "00011000",   --     **   
2373=> "00011000",   --     **   
2374=> "00011000",   --     **   
2375=> "00011000",   --     **   
-- 0xC6 ''         
2376=> "00000000",   --          
2377=> "00000000",   --          
2378=> "00000000",   --          
2379=> "00000000",   --          
2380=> "00000000",   --          
2381=> "00011111",   --     *****
2382=> "00011000",   --     **   
2383=> "00011000",   --     **   
2384=> "00011000",   --     **   
2385=> "00011000",   --     **   
2386=> "00011000",   --     **   
2387=> "00011000",   --     **   
-- 0xC7 ''         
2388=> "00011000",   --     **   
2389=> "00011000",   --     **   
2390=> "00011000",   --     **   
2391=> "00011000",   --     **   
2392=> "00011000",   --     **   
2393=> "00011111",   --     *****
2394=> "00011000",   --     **   
2395=> "00011000",   --     **   
2396=> "00011000",   --     **   
2397=> "00011000",   --     **   
2398=> "00011000",   --     **   
2399=> "00011000",   --     **   
-- 0xC8 ''         
2400=> "00000000",   --          
2401=> "00000000",   --          
2402=> "00000000",   --          
2403=> "00000000",   --          
2404=> "00000000",   --          
2405=> "11111000",   --  *****   
2406=> "00000000",   --          
2407=> "00000000",   --          
2408=> "00000000",   --          
2409=> "00000000",   --          
2410=> "00000000",   --          
2411=> "00000000",   --          
-- 0xC9 ''         
2412=> "00011000",   --     **   
2413=> "00011000",   --     **   
2414=> "00011000",   --     **   
2415=> "00011000",   --     **   
2416=> "00011000",   --     **   
2417=> "11111000",   --  *****   
2418=> "00000000",   --          
2419=> "00000000",   --          
2420=> "00000000",   --          
2421=> "00000000",   --          
2422=> "00000000",   --          
2423=> "00000000",   --          
-- 0xCA ''         
2424=> "00000000",   --          
2425=> "00000000",   --          
2426=> "00000000",   --          
2427=> "00000000",   --          
2428=> "00000000",   --          
2429=> "11111111",   --  ********
2430=> "00000000",   --          
2431=> "00000000",   --          
2432=> "00000000",   --          
2433=> "00000000",   --          
2434=> "00000000",   --          
2435=> "00000000",   --          
-- 0xCB ''         
2436=> "00011000",   --     **   
2437=> "00011000",   --     **   
2438=> "00011000",   --     **   
2439=> "00011000",   --     **   
2440=> "00011000",   --     **   
2441=> "11111111",   --  ********
2442=> "00000000",   --          
2443=> "00000000",   --          
2444=> "00000000",   --          
2445=> "00000000",   --          
2446=> "00000000",   --          
2447=> "00000000",   --          
-- 0xC C''         
2448=> "00000000",   --          
2449=> "00000000",   --          
2450=> "00000000",   --          
2451=> "00000000",   --          
2452=> "00000000",   --          
2453=> "11111000",   --  *****   
2454=> "00011000",   --     **   
2455=> "00011000",   --     **   
2456=> "00011000",   --     **   
2457=> "00011000",   --     **   
2458=> "00011000",   --     **   
2459=> "00011000",   --     **   
-- 0xCD ''         
2460=> "00011000",   --     **   
2461=> "00011000",   --     **   
2462=> "00011000",   --     **   
2463=> "00011000",   --     **   
2464=> "00011000",   --     **   
2465=> "11111000",   --  *****   
2466=> "00011000",   --     **   
2467=> "00011000",   --     **   
2468=> "00011000",   --     **   
2469=> "00011000",   --     **   
2470=> "00011000",   --     **   
2471=> "00011000",   --     **   
-- 0xCE ''         
2472=> "00000000",   --          
2473=> "00000000",   --          
2474=> "00000000",   --          
2475=> "00000000",   --          
2476=> "00000000",   --          
2477=> "11111111",   --  ********
2478=> "00011000",   --     **   
2479=> "00011000",   --     **   
2480=> "00011000",   --     **   
2481=> "00011000",   --     **   
2482=> "00011000",   --     **   
2483=> "00011000",   --     **   
-- 0xCF ''         
2484=> "00011000",   --     **   
2485=> "00011000",   --     **   
2486=> "00011000",   --     **   
2487=> "00011000",   --     **   
2488=> "00011000",   --     **   
2489=> "11111111",   --  ********
2490=> "00011000",   --     **   
2491=> "00011000",   --     **   
2492=> "00011000",   --     **   
2493=> "00011000",   --     **   
2494=> "00011000",   --     **   
2495=> "00011000",   --     **   
-- 0xD0 ''         
2496=> "00000000",   --          
2497=> "00000000",   --          
2498=> "00000000",   --          
2499=> "00000000",   --          
2500=> "00000000",   --          
2501=> "00000000",   --          
2502=> "00000000",   --          
2503=> "11111111",   --  ********
2504=> "00000000",   --          
2505=> "00000000",   --          
2506=> "00000000",   --          
2507=> "00000000",   --          
-- 0xD1 ''         
2508=> "01101100",   --   ** **  
2509=> "01101100",   --   ** **  
2510=> "01101100",   --   ** **  
2511=> "01101100",   --   ** **  
2512=> "01101100",   --   ** **  
2513=> "01101100",   --   ** **  
2514=> "01111100",   --   *****  
2515=> "00000000",   --          
2516=> "00000000",   --          
2517=> "00000000",   --          
2518=> "00000000",   --          
2519=> "00000000",   --          
-- 0xD2 ''         
2520=> "00000000",   --          
2521=> "00000000",   --          
2522=> "00000000",   --          
2523=> "00000000",   --          
2524=> "00111111",   --    ******
2525=> "00110000",   --    **    
2526=> "00111111",   --    ******
2527=> "00000000",   --          
2528=> "00000000",   --          
2529=> "00000000",   --          
2530=> "00000000",   --          
2531=> "00000000",   --          
-- 0xD3 ''         
2532=> "01101100",   --   ** **  
2533=> "01101100",   --   ** **  
2534=> "01101100",   --   ** **  
2535=> "01101100",   --   ** **  
2536=> "01101111",   --   ** ****
2537=> "01100000",   --   **     
2538=> "01111111",   --   *******
2539=> "00000000",   --          
2540=> "00000000",   --          
2541=> "00000000",   --          
2542=> "00000000",   --          
2543=> "00000000",   --          
-- 0xD4 ''         
2544=> "00000000",   --          
2545=> "00000000",   --          
2546=> "00000000",   --          
2547=> "00000000",   --          
2548=> "01111100",   --   *****  
2549=> "01101100",   --   ** **  
2550=> "01101100",   --   ** **  
2551=> "01101100",   --   ** **  
2552=> "01101100",   --   ** **  
2553=> "01101100",   --   ** **  
2554=> "01101100",   --   ** **  
2555=> "01101100",   --   ** **  
-- 0xD5 ''         
2556=> "01101100",   --   ** **  
2557=> "01101100",   --   ** **  
2558=> "01101100",   --   ** **  
2559=> "01101100",   --   ** **  
2560=> "01101100",   --   ** **  
2561=> "01101100",   --   ** **  
2562=> "01101100",   --   ** **  
2563=> "01101100",   --   ** **  
2564=> "01101100",   --   ** **  
2565=> "01101100",   --   ** **  
2566=> "01101100",   --   ** **  
2567=> "01101100",   --   ** **  
-- 0xD6 ''         
2568=> "00000000",   --          
2569=> "00000000",   --          
2570=> "00000000",   --          
2571=> "00000000",   --          
2572=> "01111111",   --   *******
2573=> "01100000",   --   **     
2574=> "01101111",   --   ** ****
2575=> "01101100",   --   ** **  
2576=> "01101100",   --   ** **  
2577=> "01101100",   --   ** **  
2578=> "01101100",   --   ** **  
2579=> "01101100",   --   ** **  
-- 0xD7 ''         
2580=> "01101100",   --   ** **  
2581=> "01101100",   --   ** **  
2582=> "01101100",   --   ** **  
2583=> "01101100",   --   ** **  
2584=> "01101111",   --   ** ****
2585=> "01100000",   --   **     
2586=> "01101111",   --   ** ****
2587=> "01101100",   --   ** **  
2588=> "01101100",   --   ** **  
2589=> "01101100",   --   ** **  
2590=> "01101100",   --   ** **  
2591=> "01101100",   --   ** **  
-- 0xD8 ''         
2592=> "00000000",   --          
2593=> "00000000",   --          
2594=> "00000000",   --          
2595=> "00000000",   --          
2596=> "11111100",   --  ******  
2597=> "00001100",   --      **  
2598=> "11111100",   --  ******  
2599=> "00000000",   --          
2600=> "00000000",   --          
2601=> "00000000",   --          
2602=> "00000000",   --          
2603=> "00000000",   --          
-- 0xD9 ''         
2604=> "01101100",   --   ** **  
2605=> "01101100",   --   ** **  
2606=> "01101100",   --   ** **  
2607=> "01101100",   --   ** **  
2608=> "11101100",   --  *** **  
2609=> "00001100",   --      **  
2610=> "11111100",   --  ******  
2611=> "00000000",   --          
2612=> "00000000",   --          
2613=> "00000000",   --          
2614=> "00000000",   --          
2615=> "00000000",   --          
-- 0xDA ''         
2616=> "00000000",   --          
2617=> "00000000",   --          
2618=> "00000000",   --          
2619=> "00000000",   --          
2620=> "11111111",   --  ********
2621=> "00000000",   --          
2622=> "11111111",   --  ********
2623=> "00000000",   --          
2624=> "00000000",   --          
2625=> "00000000",   --          
2626=> "00000000",   --          
2627=> "00000000",   --          
-- 0xDB ''         
2628=> "01101100",   --   ** **  
2629=> "01101100",   --   ** **  
2630=> "01101100",   --   ** **  
2631=> "01101100",   --   ** **  
2632=> "11101111",   --  *** ****
2633=> "00000000",   --          
2634=> "11111111",   --  ********
2635=> "00000000",   --          
2636=> "00000000",   --          
2637=> "00000000",   --          
2638=> "00000000",   --          
2639=> "00000000",   --          
-- 0xD C''         
2640=> "00000000",   --          
2641=> "00000000",   --          
2642=> "00000000",   --          
2643=> "00000000",   --          
2644=> "11111100",   --  ******  
2645=> "00001100",   --      **  
2646=> "11101100",   --  *** **  
2647=> "01101100",   --   ** **  
2648=> "01101100",   --   ** **  
2649=> "01101100",   --   ** **  
2650=> "01101100",   --   ** **  
2651=> "01101100",   --   ** **  
-- 0xDD ''         
2652=> "01101100",   --   ** **  
2653=> "01101100",   --   ** **  
2654=> "01101100",   --   ** **  
2655=> "01101100",   --   ** **  
2656=> "11101100",   --  *** **  
2657=> "00001100",   --      **  
2658=> "11101100",   --  *** **  
2659=> "01101100",   --   ** **  
2660=> "01101100",   --   ** **  
2661=> "01101100",   --   ** **  
2662=> "01101100",   --   ** **  
2663=> "01101100",   --   ** **  
-- 0xDE ''         
2664=> "00000000",   --          
2665=> "00000000",   --          
2666=> "00000000",   --          
2667=> "00000000",   --          
2668=> "11111111",   --  ********
2669=> "00000000",   --          
2670=> "11101111",   --  *** ****
2671=> "01101100",   --   ** **  
2672=> "01101100",   --   ** **  
2673=> "01101100",   --   ** **  
2674=> "01101100",   --   ** **  
2675=> "01101100",   --   ** **  
-- 0xDF ''         
2676=> "01101100",   --   ** **  
2677=> "01101100",   --   ** **  
2678=> "01101100",   --   ** **  
2679=> "01101100",   --   ** **  
2680=> "11101111",   --  *** ****
2681=> "00000000",   --          
2682=> "11101111",   --  *** ****
2683=> "01101100",   --   ** **  
2684=> "01101100",   --   ** **  
2685=> "01101100",   --   ** **  
2686=> "01101100",   --   ** **  
2687=> "01101100",   --   ** **  
-- 0xE0 ''         
2688=> "01100000",   --   **     
2689=> "00110000",   --    **    
2690=> "00011000",   --     **   
2691=> "00000000",   --          
2692=> "01111000",   --   ****   
2693=> "00001100",   --      **  
2694=> "01111100",   --   *****  
2695=> "11001100",   --  **  **  
2696=> "11011100",   --  ** ***  
2697=> "01110110",   --   *** ** 
2698=> "00000000",   --          
2699=> "00000000",   --          
-- 0xE1 ''         
2700=> "00011000",   --     **   
2701=> "00110000",   --    **    
2702=> "01100000",   --   **     
2703=> "00000000",   --          
2704=> "01111000",   --   ****   
2705=> "00001100",   --      **  
2706=> "01111100",   --   *****  
2707=> "11001100",   --  **  **  
2708=> "11011100",   --  ** ***  
2709=> "01110110",   --   *** ** 
2710=> "00000000",   --          
2711=> "00000000",   --          
-- 0xE2 ''         
2712=> "00110000",   --    **    
2713=> "01111000",   --   ****   
2714=> "11001100",   --  **  **  
2715=> "00000000",   --          
2716=> "01111000",   --   ****   
2717=> "00001100",   --      **  
2718=> "01111100",   --   *****  
2719=> "11001100",   --  **  **  
2720=> "11011100",   --  ** ***  
2721=> "01110110",   --   *** ** 
2722=> "00000000",   --          
2723=> "00000000",   --          
-- 0xE3 ''         
2724=> "00000000",   --          
2725=> "01110110",   --   *** ** 
2726=> "11011100",   --  ** ***  
2727=> "00000000",   --          
2728=> "01111000",   --   ****   
2729=> "00001100",   --      **  
2730=> "01111100",   --   *****  
2731=> "11001100",   --  **  **  
2732=> "11011100",   --  ** ***  
2733=> "01110110",   --   *** ** 
2734=> "00000000",   --          
2735=> "00000000",   --          
-- 0xE4 ''         
2736=> "00000000",   --          
2737=> "01101100",   --   ** **  
2738=> "01101100",   --   ** **  
2739=> "00000000",   --          
2740=> "01111000",   --   ****   
2741=> "00001100",   --      **  
2742=> "01111100",   --   *****  
2743=> "11001100",   --  **  **  
2744=> "11011100",   --  ** ***  
2745=> "01110110",   --   *** ** 
2746=> "00000000",   --          
2747=> "00000000",   --          
-- 0xE5 ''         
2748=> "00111000",   --    ***   
2749=> "01101100",   --   ** **  
2750=> "00111000",   --    ***   
2751=> "00000000",   --          
2752=> "01111000",   --   ****   
2753=> "00001100",   --      **  
2754=> "01111100",   --   *****  
2755=> "11001100",   --  **  **  
2756=> "11011100",   --  ** ***  
2757=> "01110110",   --   *** ** 
2758=> "00000000",   --          
2759=> "00000000",   --          
-- 0xE6 ''         
2760=> "00000000",   --          
2761=> "00000000",   --          
2762=> "00000000",   --          
2763=> "01111110",   --   ****** 
2764=> "11011011",   --  ** ** **
2765=> "00011011",   --     ** **
2766=> "01111111",   --   *******
2767=> "11011000",   --  ** **   
2768=> "11011011",   --  ** ** **
2769=> "01111110",   --   ****** 
2770=> "00000000",   --          
2771=> "00000000",   --          
-- 0xE7 ''         
2772=> "00000000",   --          
2773=> "00000000",   --          
2774=> "00000000",   --          
2775=> "01111100",   --   *****  
2776=> "11000110",   --  **   ** 
2777=> "11000000",   --  **      
2778=> "11000000",   --  **      
2779=> "11000110",   --  **   ** 
2780=> "01111100",   --   *****  
2781=> "00011000",   --     **   
2782=> "01101100",   --   ** **  
2783=> "00111000",   --    ***   
-- 0xE8 ''         
2784=> "00110000",   --    **    
2785=> "00011000",   --     **   
2786=> "00001100",   --      **  
2787=> "00000000",   --          
2788=> "01111100",   --   *****  
2789=> "11000110",   --  **   ** 
2790=> "11111110",   --  ******* 
2791=> "11000000",   --  **      
2792=> "11000110",   --  **   ** 
2793=> "01111100",   --   *****  
2794=> "00000000",   --          
2795=> "00000000",   --          
-- 0xE9 ''         
2796=> "00001100",   --      **  
2797=> "00011000",   --     **   
2798=> "00110000",   --    **    
2799=> "00000000",   --          
2800=> "01111100",   --   *****  
2801=> "11000110",   --  **   ** 
2802=> "11111110",   --  ******* 
2803=> "11000000",   --  **      
2804=> "11000110",   --  **   ** 
2805=> "01111100",   --   *****  
2806=> "00000000",   --          
2807=> "00000000",   --          
-- 0xEA ''         
2808=> "00010000",   --     *    
2809=> "00111000",   --    ***   
2810=> "01101100",   --   ** **  
2811=> "00000000",   --          
2812=> "01111100",   --   *****  
2813=> "11000110",   --  **   ** 
2814=> "11111110",   --  ******* 
2815=> "11000000",   --  **      
2816=> "11000110",   --  **   ** 
2817=> "01111100",   --   *****  
2818=> "00000000",   --          
2819=> "00000000",   --          
-- 0xEB ''         
2820=> "00000000",   --          
2821=> "01101100",   --   ** **  
2822=> "01101100",   --   ** **  
2823=> "00000000",   --          
2824=> "01111100",   --   *****  
2825=> "11000110",   --  **   ** 
2826=> "11111110",   --  ******* 
2827=> "11000000",   --  **      
2828=> "11000110",   --  **   ** 
2829=> "01111100",   --   *****  
2830=> "00000000",   --          
2831=> "00000000",   --          
-- 0xE C''         
2832=> "01100000",   --   **     
2833=> "00110000",   --    **    
2834=> "00011000",   --     **   
2835=> "00000000",   --          
2836=> "00111000",   --    ***   
2837=> "00011000",   --     **   
2838=> "00011000",   --     **   
2839=> "00011000",   --     **   
2840=> "00011000",   --     **   
2841=> "00111100",   --    ****  
2842=> "00000000",   --          
2843=> "00000000",   --          
-- 0xED ''         
2844=> "00001100",   --      **  
2845=> "00011000",   --     **   
2846=> "00110000",   --    **    
2847=> "00000000",   --          
2848=> "00111000",   --    ***   
2849=> "00011000",   --     **   
2850=> "00011000",   --     **   
2851=> "00011000",   --     **   
2852=> "00011000",   --     **   
2853=> "00111100",   --    ****  
2854=> "00000000",   --          
2855=> "00000000",   --          
-- 0xEE ''         
2856=> "00011000",   --     **   
2857=> "00111100",   --    ****  
2858=> "01100110",   --   **  ** 
2859=> "00000000",   --          
2860=> "00111000",   --    ***   
2861=> "00011000",   --     **   
2862=> "00011000",   --     **   
2863=> "00011000",   --     **   
2864=> "00011000",   --     **   
2865=> "00111100",   --    ****  
2866=> "00000000",   --          
2867=> "00000000",   --          
-- 0xEF ''         
2868=> "00000000",   --          
2869=> "01101100",   --   ** **  
2870=> "01101100",   --   ** **  
2871=> "00000000",   --          
2872=> "00111000",   --    ***   
2873=> "00011000",   --     **   
2874=> "00011000",   --     **   
2875=> "00011000",   --     **   
2876=> "00011000",   --     **   
2877=> "00111100",   --    ****  
2878=> "00000000",   --          
2879=> "00000000",   --          
-- 0xF0 ''         
2880=> "01111000",   --   ****   
2881=> "00110000",   --    **    
2882=> "01111000",   --   ****   
2883=> "00001100",   --      **  
2884=> "01111110",   --   ****** 
2885=> "11000110",   --  **   ** 
2886=> "11000110",   --  **   ** 
2887=> "11000110",   --  **   ** 
2888=> "11000110",   --  **   ** 
2889=> "01111100",   --   *****  
2890=> "00000000",   --          
2891=> "00000000",   --          
-- 0xF1 ''         
2892=> "00000000",   --          
2893=> "01110110",   --   *** ** 
2894=> "11011100",   --  ** ***  
2895=> "00000000",   --          
2896=> "11011100",   --  ** ***  
2897=> "01100110",   --   **  ** 
2898=> "01100110",   --   **  ** 
2899=> "01100110",   --   **  ** 
2900=> "01100110",   --   **  ** 
2901=> "01100110",   --   **  ** 
2902=> "00000000",   --          
2903=> "00000000",   --          
-- 0xF2 ''         
2904=> "01100000",   --   **     
2905=> "00110000",   --    **    
2906=> "00011000",   --     **   
2907=> "00000000",   --          
2908=> "01111100",   --   *****  
2909=> "11000110",   --  **   ** 
2910=> "11000110",   --  **   ** 
2911=> "11000110",   --  **   ** 
2912=> "11000110",   --  **   ** 
2913=> "01111100",   --   *****  
2914=> "00000000",   --          
2915=> "00000000",   --          
-- 0xF3 ''         
2916=> "00001100",   --      **  
2917=> "00011000",   --     **   
2918=> "00110000",   --    **    
2919=> "00000000",   --          
2920=> "01111100",   --   *****  
2921=> "11000110",   --  **   ** 
2922=> "11000110",   --  **   ** 
2923=> "11000110",   --  **   ** 
2924=> "11000110",   --  **   ** 
2925=> "01111100",   --   *****  
2926=> "00000000",   --          
2927=> "00000000",   --          
-- 0xF4 ''         
2928=> "00010000",   --     *    
2929=> "00111000",   --    ***   
2930=> "01101100",   --   ** **  
2931=> "00000000",   --          
2932=> "01111100",   --   *****  
2933=> "11000110",   --  **   ** 
2934=> "11000110",   --  **   ** 
2935=> "11000110",   --  **   ** 
2936=> "11000110",   --  **   ** 
2937=> "01111100",   --   *****  
2938=> "00000000",   --          
2939=> "00000000",   --          
-- 0xF5 ''         
2940=> "00000000",   --          
2941=> "01110110",   --   *** ** 
2942=> "11011100",   --  ** ***  
2943=> "00000000",   --          
2944=> "01111100",   --   *****  
2945=> "11000110",   --  **   ** 
2946=> "11000110",   --  **   ** 
2947=> "11000110",   --  **   ** 
2948=> "11000110",   --  **   ** 
2949=> "01111100",   --   *****  
2950=> "00000000",   --          
2951=> "00000000",   --          
-- 0xF6 ''         
2952=> "00000000",   --          
2953=> "01101100",   --   ** **  
2954=> "01101100",   --   ** **  
2955=> "00000000",   --          
2956=> "01111100",   --   *****  
2957=> "11000110",   --  **   ** 
2958=> "11000110",   --  **   ** 
2959=> "11000110",   --  **   ** 
2960=> "11000110",   --  **   ** 
2961=> "01111100",   --   *****  
2962=> "00000000",   --          
2963=> "00000000",   --          
-- 0xF7 ''         
2964=> "00000000",   --          
2965=> "00000000",   --          
2966=> "00011000",   --     **   
2967=> "00011000",   --     **   
2968=> "00000000",   --          
2969=> "01111110",   --   ****** 
2970=> "00000000",   --          
2971=> "00011000",   --     **   
2972=> "00011000",   --     **   
2973=> "00000000",   --          
2974=> "00000000",   --          
2975=> "00000000",   --          
-- 0xF8 ''         
2976=> "00000000",   --          
2977=> "00000000",   --          
2978=> "00000000",   --          
2979=> "00000000",   --          
2980=> "01111110",   --   ****** 
2981=> "11001110",   --  **  *** 
2982=> "11011110",   --  ** **** 
2983=> "11110110",   --  **** ** 
2984=> "11100110",   --  ***  ** 
2985=> "11111100",   --  ******  
2986=> "00000000",   --          
2987=> "00000000",   --          
-- 0xF9 ''         
2988=> "11000000",   --  **      
2989=> "01100000",   --   **     
2990=> "00110000",   --    **    
2991=> "00000000",   --          
2992=> "11001100",   --  **  **  
2993=> "11001100",   --  **  **  
2994=> "11001100",   --  **  **  
2995=> "11001100",   --  **  **  
2996=> "11001100",   --  **  **  
2997=> "01110110",   --   *** ** 
2998=> "00000000",   --          
2999=> "00000000",   --          
-- 0xFA ''         
3000=> "00001100",   --      **  
3001=> "00011000",   --     **   
3002=> "00110000",   --    **    
3003=> "00000000",   --          
3004=> "11001100",   --  **  **  
3005=> "11001100",   --  **  **  
3006=> "11001100",   --  **  **  
3007=> "11001100",   --  **  **  
3008=> "11001100",   --  **  **  
3009=> "01110110",   --   *** ** 
3010=> "00000000",   --          
3011=> "00000000",   --          
-- 0xFB ''         
3012=> "00110000",   --    **    
3013=> "01111000",   --   ****   
3014=> "11001100",   --  **  **  
3015=> "00000000",   --          
3016=> "11001100",   --  **  **  
3017=> "11001100",   --  **  **  
3018=> "11001100",   --  **  **  
3019=> "11001100",   --  **  **  
3020=> "11001100",   --  **  **  
3021=> "01110110",   --   *** ** 
3022=> "00000000",   --          
3023=> "00000000",   --          
-- 0xFC ''         
3024=> "00000000",   --          
3025=> "11001100",   --  **  **  
3026=> "11001100",   --  **  **  
3027=> "00000000",   --          
3028=> "11001100",   --  **  **  
3029=> "11001100",   --  **  **  
3030=> "11001100",   --  **  **  
3031=> "11001100",   --  **  **  
3032=> "11001100",   --  **  **  
3033=> "01110110",   --   *** ** 
3034=> "00000000",   --          
3035=> "00000000",   --          
-- 0xFD ''         
3036=> "00001100",   --      **  
3037=> "00011000",   --     **   
3038=> "00110000",   --    **    
3039=> "00000000",   --          
3040=> "11000110",   --  **   ** 
3041=> "11000110",   --  **   ** 
3042=> "11000110",   --  **   ** 
3043=> "11001110",   --  **  *** 
3044=> "01110110",   --   *** ** 
3045=> "00000110",   --       ** 
3046=> "11000110",   --  **   ** 
3047=> "01111100",   --   *****  
-- 0xFE ''         
3048=> "00000000",   --          
3049=> "11110000",   --  ****    
3050=> "01100000",   --   **     
3051=> "01100000",   --   **     
3052=> "01111000",   --   ****   
3053=> "01101100",   --   ** **  
3054=> "01101100",   --   ** **  
3055=> "01101100",   --   ** **  
3056=> "01111000",   --   ****   
3057=> "01100000",   --   **     
3058=> "01100000",   --   **     
3059=> "11110000",   --  ****    
-- 0xFF ''         
3060=> "00000000",   --          
3061=> "11000110",   --  **   ** 
3062=> "11000110",   --  **   ** 
3063=> "00000000",   --          
3064=> "11000110",   --  **   ** 
3065=> "11000110",   --  **   ** 
3066=> "11000110",   --  **   ** 
3067=> "11001110",   --  **  *** 
3068=> "01110110",   --   *** ** 
3069=> "00000110",   --       ** 
3070=> "11000110",   --  **   ** 
3071=> "01111100",   --   *****  
--
others => "00000000"
);


begin
    rom : process (clk)
    begin
        if rising_edge(clk) then
            data_out <=mem(to_integer(unsigned(address)));
        end if;
    end process rom;

    --data_out <=mem(to_integer(unsigned(address)));

end architecture synth;